// This is the unpowered netlist.
module simd (clk,
    data_R,
    data_W,
    done,
    rst,
    data_address,
    data_in,
    data_out,
    instruction_address,
    instruction_in);
 input clk;
 output data_R;
 output data_W;
 output done;
 input rst;
 output [9:0] data_address;
 input [15:0] data_in;
 output [15:0] data_out;
 output [9:0] instruction_address;
 input [17:0] instruction_in;

 wire \Add.sub ;
 wire CMD_addition;
 wire CMD_and;
 wire CMD_load;
 wire CMD_logic_shift_right;
 wire CMD_loopjump;
 wire CMD_mul_accumulation;
 wire CMD_multiplication;
 wire CMD_not;
 wire CMD_or;
 wire CMD_set;
 wire CMD_setloop;
 wire CMD_store;
 wire \H[0][0] ;
 wire \H[0][10] ;
 wire \H[0][11] ;
 wire \H[0][12] ;
 wire \H[0][13] ;
 wire \H[0][14] ;
 wire \H[0][15] ;
 wire \H[0][1] ;
 wire \H[0][2] ;
 wire \H[0][3] ;
 wire \H[0][4] ;
 wire \H[0][5] ;
 wire \H[0][6] ;
 wire \H[0][7] ;
 wire \H[0][8] ;
 wire \H[0][9] ;
 wire \H[1][0] ;
 wire \H[1][10] ;
 wire \H[1][11] ;
 wire \H[1][12] ;
 wire \H[1][13] ;
 wire \H[1][14] ;
 wire \H[1][15] ;
 wire \H[1][1] ;
 wire \H[1][2] ;
 wire \H[1][3] ;
 wire \H[1][4] ;
 wire \H[1][5] ;
 wire \H[1][6] ;
 wire \H[1][7] ;
 wire \H[1][8] ;
 wire \H[1][9] ;
 wire \H[2][0] ;
 wire \H[2][10] ;
 wire \H[2][11] ;
 wire \H[2][12] ;
 wire \H[2][13] ;
 wire \H[2][14] ;
 wire \H[2][15] ;
 wire \H[2][1] ;
 wire \H[2][2] ;
 wire \H[2][3] ;
 wire \H[2][4] ;
 wire \H[2][5] ;
 wire \H[2][6] ;
 wire \H[2][7] ;
 wire \H[2][8] ;
 wire \H[2][9] ;
 wire \H[3][0] ;
 wire \H[3][10] ;
 wire \H[3][11] ;
 wire \H[3][12] ;
 wire \H[3][13] ;
 wire \H[3][14] ;
 wire \H[3][15] ;
 wire \H[3][1] ;
 wire \H[3][2] ;
 wire \H[3][3] ;
 wire \H[3][4] ;
 wire \H[3][5] ;
 wire \H[3][6] ;
 wire \H[3][7] ;
 wire \H[3][8] ;
 wire \H[3][9] ;
 wire Him;
 wire Hreg2;
 wire Hreg3;
 wire \LC[0] ;
 wire \LC[1] ;
 wire \LC[2] ;
 wire \LC[3] ;
 wire \LC[4] ;
 wire \LC[5] ;
 wire \LC[6] ;
 wire \LC[7] ;
 wire \LC[8] ;
 wire \LC[9] ;
 wire Oim;
 wire Oreg2;
 wire Oreg3;
 wire \Oset[0][0] ;
 wire \Oset[0][10] ;
 wire \Oset[0][11] ;
 wire \Oset[0][12] ;
 wire \Oset[0][13] ;
 wire \Oset[0][14] ;
 wire \Oset[0][15] ;
 wire \Oset[0][1] ;
 wire \Oset[0][2] ;
 wire \Oset[0][3] ;
 wire \Oset[0][4] ;
 wire \Oset[0][5] ;
 wire \Oset[0][6] ;
 wire \Oset[0][7] ;
 wire \Oset[0][8] ;
 wire \Oset[0][9] ;
 wire \Oset[1][0] ;
 wire \Oset[1][10] ;
 wire \Oset[1][11] ;
 wire \Oset[1][12] ;
 wire \Oset[1][13] ;
 wire \Oset[1][14] ;
 wire \Oset[1][15] ;
 wire \Oset[1][1] ;
 wire \Oset[1][2] ;
 wire \Oset[1][3] ;
 wire \Oset[1][4] ;
 wire \Oset[1][5] ;
 wire \Oset[1][6] ;
 wire \Oset[1][7] ;
 wire \Oset[1][8] ;
 wire \Oset[1][9] ;
 wire \Oset[2][0] ;
 wire \Oset[2][10] ;
 wire \Oset[2][11] ;
 wire \Oset[2][12] ;
 wire \Oset[2][13] ;
 wire \Oset[2][14] ;
 wire \Oset[2][15] ;
 wire \Oset[2][1] ;
 wire \Oset[2][2] ;
 wire \Oset[2][3] ;
 wire \Oset[2][4] ;
 wire \Oset[2][5] ;
 wire \Oset[2][6] ;
 wire \Oset[2][7] ;
 wire \Oset[2][8] ;
 wire \Oset[2][9] ;
 wire \Oset[3][0] ;
 wire \Oset[3][10] ;
 wire \Oset[3][11] ;
 wire \Oset[3][12] ;
 wire \Oset[3][13] ;
 wire \Oset[3][14] ;
 wire \Oset[3][15] ;
 wire \Oset[3][1] ;
 wire \Oset[3][2] ;
 wire \Oset[3][3] ;
 wire \Oset[3][4] ;
 wire \Oset[3][5] ;
 wire \Oset[3][6] ;
 wire \Oset[3][7] ;
 wire \Oset[3][8] ;
 wire \Oset[3][9] ;
 wire Qim;
 wire Qreg2;
 wire Qreg3;
 wire \Qset[0][0] ;
 wire \Qset[0][10] ;
 wire \Qset[0][11] ;
 wire \Qset[0][12] ;
 wire \Qset[0][13] ;
 wire \Qset[0][14] ;
 wire \Qset[0][15] ;
 wire \Qset[0][1] ;
 wire \Qset[0][2] ;
 wire \Qset[0][3] ;
 wire \Qset[0][4] ;
 wire \Qset[0][5] ;
 wire \Qset[0][6] ;
 wire \Qset[0][7] ;
 wire \Qset[0][8] ;
 wire \Qset[0][9] ;
 wire \Qset[1][0] ;
 wire \Qset[1][10] ;
 wire \Qset[1][11] ;
 wire \Qset[1][12] ;
 wire \Qset[1][13] ;
 wire \Qset[1][14] ;
 wire \Qset[1][15] ;
 wire \Qset[1][1] ;
 wire \Qset[1][2] ;
 wire \Qset[1][3] ;
 wire \Qset[1][4] ;
 wire \Qset[1][5] ;
 wire \Qset[1][6] ;
 wire \Qset[1][7] ;
 wire \Qset[1][8] ;
 wire \Qset[1][9] ;
 wire \Qset[2][0] ;
 wire \Qset[2][10] ;
 wire \Qset[2][11] ;
 wire \Qset[2][12] ;
 wire \Qset[2][13] ;
 wire \Qset[2][14] ;
 wire \Qset[2][15] ;
 wire \Qset[2][1] ;
 wire \Qset[2][2] ;
 wire \Qset[2][3] ;
 wire \Qset[2][4] ;
 wire \Qset[2][5] ;
 wire \Qset[2][6] ;
 wire \Qset[2][7] ;
 wire \Qset[2][8] ;
 wire \Qset[2][9] ;
 wire \Qset[3][0] ;
 wire \Qset[3][10] ;
 wire \Qset[3][11] ;
 wire \Qset[3][12] ;
 wire \Qset[3][13] ;
 wire \Qset[3][14] ;
 wire \Qset[3][15] ;
 wire \Qset[3][1] ;
 wire \Qset[3][2] ;
 wire \Qset[3][3] ;
 wire \Qset[3][4] ;
 wire \Qset[3][5] ;
 wire \Qset[3][6] ;
 wire \Qset[3][7] ;
 wire \Qset[3][8] ;
 wire \Qset[3][9] ;
 wire \R0[0] ;
 wire \R0[1] ;
 wire \R1[0] ;
 wire \R1[1] ;
 wire \R2[0] ;
 wire \R2[1] ;
 wire \R3[0] ;
 wire \R3[1] ;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire \current_state[0] ;
 wire \current_state[1] ;
 wire \current_state[2] ;
 wire \current_state[4] ;
 wire \current_state[5] ;
 wire \current_state[6] ;
 wire \im_reg[6] ;
 wire \im_reg[7] ;
 wire \im_reg[8] ;
 wire \im_reg[9] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net8;
 wire net9;
 wire \next_PC[0] ;
 wire \next_PC[1] ;
 wire \next_PC[2] ;
 wire \next_PC[3] ;
 wire \next_PC[4] ;
 wire \next_PC[5] ;
 wire \next_PC[6] ;
 wire \next_PC[7] ;
 wire \next_PC[8] ;
 wire \next_PC[9] ;
 wire \result_reg_Lshift[0] ;
 wire \result_reg_Lshift[10] ;
 wire \result_reg_Lshift[11] ;
 wire \result_reg_Lshift[12] ;
 wire \result_reg_Lshift[13] ;
 wire \result_reg_Lshift[14] ;
 wire \result_reg_Lshift[15] ;
 wire \result_reg_Lshift[1] ;
 wire \result_reg_Lshift[2] ;
 wire \result_reg_Lshift[3] ;
 wire \result_reg_Lshift[4] ;
 wire \result_reg_Lshift[5] ;
 wire \result_reg_Lshift[6] ;
 wire \result_reg_Lshift[7] ;
 wire \result_reg_Lshift[8] ;
 wire \result_reg_Lshift[9] ;
 wire \result_reg_Rshift[0] ;
 wire \result_reg_Rshift[10] ;
 wire \result_reg_Rshift[11] ;
 wire \result_reg_Rshift[12] ;
 wire \result_reg_Rshift[13] ;
 wire \result_reg_Rshift[14] ;
 wire \result_reg_Rshift[15] ;
 wire \result_reg_Rshift[1] ;
 wire \result_reg_Rshift[2] ;
 wire \result_reg_Rshift[3] ;
 wire \result_reg_Rshift[4] ;
 wire \result_reg_Rshift[5] ;
 wire \result_reg_Rshift[6] ;
 wire \result_reg_Rshift[7] ;
 wire \result_reg_Rshift[8] ;
 wire \result_reg_Rshift[9] ;
 wire \result_reg_add[0] ;
 wire \result_reg_add[10] ;
 wire \result_reg_add[11] ;
 wire \result_reg_add[12] ;
 wire \result_reg_add[13] ;
 wire \result_reg_add[14] ;
 wire \result_reg_add[15] ;
 wire \result_reg_add[1] ;
 wire \result_reg_add[2] ;
 wire \result_reg_add[3] ;
 wire \result_reg_add[4] ;
 wire \result_reg_add[5] ;
 wire \result_reg_add[6] ;
 wire \result_reg_add[7] ;
 wire \result_reg_add[8] ;
 wire \result_reg_add[9] ;
 wire \result_reg_and[0] ;
 wire \result_reg_and[10] ;
 wire \result_reg_and[11] ;
 wire \result_reg_and[12] ;
 wire \result_reg_and[13] ;
 wire \result_reg_and[14] ;
 wire \result_reg_and[15] ;
 wire \result_reg_and[1] ;
 wire \result_reg_and[2] ;
 wire \result_reg_and[3] ;
 wire \result_reg_and[4] ;
 wire \result_reg_and[5] ;
 wire \result_reg_and[6] ;
 wire \result_reg_and[7] ;
 wire \result_reg_and[8] ;
 wire \result_reg_and[9] ;
 wire \result_reg_mac[0] ;
 wire \result_reg_mac[10] ;
 wire \result_reg_mac[11] ;
 wire \result_reg_mac[12] ;
 wire \result_reg_mac[13] ;
 wire \result_reg_mac[14] ;
 wire \result_reg_mac[15] ;
 wire \result_reg_mac[1] ;
 wire \result_reg_mac[2] ;
 wire \result_reg_mac[3] ;
 wire \result_reg_mac[4] ;
 wire \result_reg_mac[5] ;
 wire \result_reg_mac[6] ;
 wire \result_reg_mac[7] ;
 wire \result_reg_mac[8] ;
 wire \result_reg_mac[9] ;
 wire \result_reg_mul[0] ;
 wire \result_reg_mul[10] ;
 wire \result_reg_mul[11] ;
 wire \result_reg_mul[12] ;
 wire \result_reg_mul[13] ;
 wire \result_reg_mul[14] ;
 wire \result_reg_mul[15] ;
 wire \result_reg_mul[1] ;
 wire \result_reg_mul[2] ;
 wire \result_reg_mul[3] ;
 wire \result_reg_mul[4] ;
 wire \result_reg_mul[5] ;
 wire \result_reg_mul[6] ;
 wire \result_reg_mul[7] ;
 wire \result_reg_mul[8] ;
 wire \result_reg_mul[9] ;
 wire \result_reg_not[0] ;
 wire \result_reg_not[10] ;
 wire \result_reg_not[11] ;
 wire \result_reg_not[12] ;
 wire \result_reg_not[13] ;
 wire \result_reg_not[14] ;
 wire \result_reg_not[15] ;
 wire \result_reg_not[1] ;
 wire \result_reg_not[2] ;
 wire \result_reg_not[3] ;
 wire \result_reg_not[4] ;
 wire \result_reg_not[5] ;
 wire \result_reg_not[6] ;
 wire \result_reg_not[7] ;
 wire \result_reg_not[8] ;
 wire \result_reg_not[9] ;
 wire \result_reg_or[0] ;
 wire \result_reg_or[10] ;
 wire \result_reg_or[11] ;
 wire \result_reg_or[12] ;
 wire \result_reg_or[13] ;
 wire \result_reg_or[14] ;
 wire \result_reg_or[15] ;
 wire \result_reg_or[1] ;
 wire \result_reg_or[2] ;
 wire \result_reg_or[3] ;
 wire \result_reg_or[4] ;
 wire \result_reg_or[5] ;
 wire \result_reg_or[6] ;
 wire \result_reg_or[7] ;
 wire \result_reg_or[8] ;
 wire \result_reg_or[9] ;
 wire \result_reg_set[0] ;
 wire \result_reg_set[10] ;
 wire \result_reg_set[11] ;
 wire \result_reg_set[12] ;
 wire \result_reg_set[13] ;
 wire \result_reg_set[14] ;
 wire \result_reg_set[15] ;
 wire \result_reg_set[1] ;
 wire \result_reg_set[2] ;
 wire \result_reg_set[3] ;
 wire \result_reg_set[4] ;
 wire \result_reg_set[5] ;
 wire \result_reg_set[6] ;
 wire \result_reg_set[7] ;
 wire \result_reg_set[8] ;
 wire \result_reg_set[9] ;
 wire \result_reg_sub[0] ;
 wire \result_reg_sub[10] ;
 wire \result_reg_sub[11] ;
 wire \result_reg_sub[12] ;
 wire \result_reg_sub[13] ;
 wire \result_reg_sub[14] ;
 wire \result_reg_sub[15] ;
 wire \result_reg_sub[1] ;
 wire \result_reg_sub[2] ;
 wire \result_reg_sub[3] ;
 wire \result_reg_sub[4] ;
 wire \result_reg_sub[5] ;
 wire \result_reg_sub[6] ;
 wire \result_reg_sub[7] ;
 wire \result_reg_sub[8] ;
 wire \result_reg_sub[9] ;
 wire \shift.H ;
 wire \shift.O ;
 wire \shift.Q ;
 wire \shift.left ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_00073_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_00649_));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(_01823_));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(_01830_));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(_01834_));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(_01850_));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(_01870_));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(_01890_));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(_01909_));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(_01914_));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(_01929_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_00677_));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(_02168_));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(_02168_));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(_02382_));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(_02474_));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(_02545_));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(_02545_));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(_02840_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_00677_));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(_03449_));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(_03601_));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(_03601_));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(_04721_));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(_05115_));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(_05115_));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(_05298_));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(_05298_));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(_05693_));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(_05711_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_00683_));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(_05717_));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(_05725_));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(_06012_));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(_06030_));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(_06182_));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(_06218_));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(_06218_));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(_06218_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_00717_));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(_06218_));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(\im_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(\im_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(\im_reg[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(\result_reg_mac[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_00722_));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(\R2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(\R2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(\R2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(\R2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(\R2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(\R2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(\R2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(\R2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_00742_));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(\R2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(\R3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(\R3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(_00396_));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(_00498_));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(_00498_));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(_00997_));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(_01047_));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(_01285_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_00750_));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(_01332_));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(_01332_));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(_01362_));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(_01670_));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(_01771_));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(_01785_));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(_01883_));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(_01905_));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(_02101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_00759_));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(_03136_));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(_05634_));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(_05634_));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(\im_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(_00809_));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(_00809_));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(_00809_));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(_00809_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_00759_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_00473_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_00759_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_00776_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_00802_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_00814_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_00818_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_00820_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_00846_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_00871_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_00878_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_00498_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_00878_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_00904_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_00904_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_00904_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_00909_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_00946_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_00953_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_00953_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_00953_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_00972_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_00564_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_01044_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_01072_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_01074_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(_01085_));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_01098_));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_01149_));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_01149_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_01149_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_01150_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_00567_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_01205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_01270_));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_01278_));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(_01284_));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(_01325_));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(_01349_));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_01349_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(_01368_));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(_01368_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_00621_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_01368_));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_01380_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(_01396_));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(_01410_));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(_01437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(_01437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(_01437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(_01444_));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(_01462_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_00621_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(_01467_));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(_01485_));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(_01488_));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(_01496_));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(_01502_));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(_01507_));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(_01591_));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(_01621_));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(_01668_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_00626_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(_01690_));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(_01711_));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(_01712_));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(_01727_));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(_01731_));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(_01757_));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(_01768_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_00648_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(_01775_));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(_01788_));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(_01792_));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(_01801_));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(_01801_));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(_01806_));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(_01811_));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(_01819_));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(_01819_));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(_01819_));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_332 ();
 sky130_fd_sc_hd__inv_2 _06286_ (.A(net25),
    .Y(_06253_));
 sky130_fd_sc_hd__nand2_1 _06287_ (.A(net23),
    .B(net24),
    .Y(_06254_));
 sky130_fd_sc_hd__nand2_1 _06288_ (.A(net20),
    .B(net21),
    .Y(_06255_));
 sky130_fd_sc_hd__inv_2 _06289_ (.A(_06255_),
    .Y(_06256_));
 sky130_fd_sc_hd__nand2_1 _06290_ (.A(_06256_),
    .B(net22),
    .Y(_06257_));
 sky130_fd_sc_hd__or3_2 _06291_ (.A(_06253_),
    .B(_06254_),
    .C(_06257_),
    .X(_06258_));
 sky130_fd_sc_hd__inv_2 _06292_ (.A(net35),
    .Y(_06259_));
 sky130_fd_sc_hd__nand2_1 _06293_ (.A(_06259_),
    .B(net64),
    .Y(_06260_));
 sky130_fd_sc_hd__o21ai_1 _06294_ (.A1(net35),
    .A2(_06258_),
    .B1(_06260_),
    .Y(_00013_));
 sky130_fd_sc_hd__nand2_1 _06295_ (.A(_06258_),
    .B(_06259_),
    .Y(_06261_));
 sky130_fd_sc_hd__or2b_1 _06296_ (.A(_06261_),
    .B_N(\current_state[1] ),
    .X(_06262_));
 sky130_fd_sc_hd__inv_2 _06297_ (.A(_06262_),
    .Y(_00011_));
 sky130_fd_sc_hd__inv_2 _06298_ (.A(\current_state[0] ),
    .Y(_06263_));
 sky130_fd_sc_hd__inv_2 _06299_ (.A(\current_state[5] ),
    .Y(_06264_));
 sky130_fd_sc_hd__a21o_1 _06300_ (.A1(_06263_),
    .A2(_06264_),
    .B1(_06261_),
    .X(_06265_));
 sky130_fd_sc_hd__inv_2 _06301_ (.A(_06265_),
    .Y(_00010_));
 sky130_fd_sc_hd__inv_2 _06302_ (.A(\current_state[2] ),
    .Y(_06266_));
 sky130_fd_sc_hd__clkbuf_4 _06303_ (.A(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__or2_1 _06304_ (.A(_06267_),
    .B(_06261_),
    .X(_06268_));
 sky130_fd_sc_hd__inv_2 _06305_ (.A(_06268_),
    .Y(_00012_));
 sky130_fd_sc_hd__inv_2 _06306_ (.A(\current_state[6] ),
    .Y(_06269_));
 sky130_fd_sc_hd__or2_1 _06307_ (.A(_06269_),
    .B(_06261_),
    .X(_06270_));
 sky130_fd_sc_hd__inv_2 _06308_ (.A(_06270_),
    .Y(_00008_));
 sky130_fd_sc_hd__inv_2 _06309_ (.A(\current_state[4] ),
    .Y(_06271_));
 sky130_fd_sc_hd__or2_1 _06310_ (.A(_06271_),
    .B(_06261_),
    .X(_06272_));
 sky130_fd_sc_hd__inv_2 _06311_ (.A(_06272_),
    .Y(_00009_));
 sky130_fd_sc_hd__or2_1 _06312_ (.A(\LC[1] ),
    .B(\LC[0] ),
    .X(_06273_));
 sky130_fd_sc_hd__or2_1 _06313_ (.A(\LC[2] ),
    .B(_06273_),
    .X(_06274_));
 sky130_fd_sc_hd__or2_1 _06314_ (.A(\LC[3] ),
    .B(_06274_),
    .X(_06275_));
 sky130_fd_sc_hd__nor2_1 _06315_ (.A(\LC[4] ),
    .B(_06275_),
    .Y(_06276_));
 sky130_fd_sc_hd__inv_2 _06316_ (.A(_06276_),
    .Y(_06277_));
 sky130_fd_sc_hd__nor2_1 _06317_ (.A(\LC[5] ),
    .B(_06277_),
    .Y(_06278_));
 sky130_fd_sc_hd__inv_2 _06318_ (.A(_06278_),
    .Y(_06279_));
 sky130_fd_sc_hd__nor2_1 _06319_ (.A(\LC[6] ),
    .B(_06279_),
    .Y(_06280_));
 sky130_fd_sc_hd__and2b_1 _06320_ (.A_N(\LC[7] ),
    .B(_06280_),
    .X(_06281_));
 sky130_fd_sc_hd__inv_2 _06321_ (.A(\LC[8] ),
    .Y(_06282_));
 sky130_fd_sc_hd__nand2_2 _06322_ (.A(_06281_),
    .B(_06282_),
    .Y(_06283_));
 sky130_fd_sc_hd__o21ai_4 _06323_ (.A1(\LC[9] ),
    .A2(_06283_),
    .B1(CMD_loopjump),
    .Y(_06284_));
 sky130_fd_sc_hd__buf_2 _06324_ (.A(_06284_),
    .X(_06285_));
 sky130_fd_sc_hd__or2_1 _06325_ (.A(\R3[0] ),
    .B(_06285_),
    .X(_00470_));
 sky130_fd_sc_hd__and3_2 _06326_ (.A(_06259_),
    .B(_06263_),
    .C(_06271_),
    .X(_00471_));
 sky130_fd_sc_hd__buf_2 _06327_ (.A(_00471_),
    .X(_00472_));
 sky130_fd_sc_hd__nand2_2 _06328_ (.A(_00472_),
    .B(\current_state[6] ),
    .Y(_00473_));
 sky130_fd_sc_hd__inv_2 _06329_ (.A(_00473_),
    .Y(_00474_));
 sky130_fd_sc_hd__clkbuf_4 _06330_ (.A(_00474_),
    .X(_00475_));
 sky130_fd_sc_hd__nand2_1 _06331_ (.A(_06285_),
    .B(\next_PC[0] ),
    .Y(_00476_));
 sky130_fd_sc_hd__nand2_1 _06332_ (.A(_00473_),
    .B(_06259_),
    .Y(_00477_));
 sky130_fd_sc_hd__inv_2 _06333_ (.A(_00477_),
    .Y(_00478_));
 sky130_fd_sc_hd__a32o_1 _06334_ (.A1(_00470_),
    .A2(_00475_),
    .A3(_00476_),
    .B1(\next_PC[0] ),
    .B2(_00478_),
    .X(_00014_));
 sky130_fd_sc_hd__or2_1 _06335_ (.A(\R3[1] ),
    .B(_06285_),
    .X(_00479_));
 sky130_fd_sc_hd__nand2_1 _06336_ (.A(\next_PC[1] ),
    .B(\next_PC[0] ),
    .Y(_00480_));
 sky130_fd_sc_hd__inv_2 _06337_ (.A(_00480_),
    .Y(_00481_));
 sky130_fd_sc_hd__nor2_1 _06338_ (.A(\next_PC[1] ),
    .B(\next_PC[0] ),
    .Y(_00482_));
 sky130_fd_sc_hd__o21ai_1 _06339_ (.A1(_00481_),
    .A2(_00482_),
    .B1(_06285_),
    .Y(_00483_));
 sky130_fd_sc_hd__a32o_1 _06340_ (.A1(_00479_),
    .A2(_00475_),
    .A3(_00483_),
    .B1(\next_PC[1] ),
    .B2(_00478_),
    .X(_00015_));
 sky130_fd_sc_hd__nand2_1 _06341_ (.A(_00481_),
    .B(\next_PC[2] ),
    .Y(_00484_));
 sky130_fd_sc_hd__or2_1 _06342_ (.A(\next_PC[2] ),
    .B(_00481_),
    .X(_00485_));
 sky130_fd_sc_hd__buf_2 _06343_ (.A(_06284_),
    .X(_00486_));
 sky130_fd_sc_hd__a21bo_1 _06344_ (.A1(_00484_),
    .A2(_00485_),
    .B1_N(_00486_),
    .X(_00487_));
 sky130_fd_sc_hd__or2_1 _06345_ (.A(\R2[0] ),
    .B(_00486_),
    .X(_00488_));
 sky130_fd_sc_hd__a32o_1 _06346_ (.A1(_00487_),
    .A2(_00475_),
    .A3(_00488_),
    .B1(\next_PC[2] ),
    .B2(_00478_),
    .X(_00016_));
 sky130_fd_sc_hd__or2_1 _06347_ (.A(\R2[1] ),
    .B(_06285_),
    .X(_00489_));
 sky130_fd_sc_hd__inv_2 _06348_ (.A(\next_PC[3] ),
    .Y(_00490_));
 sky130_fd_sc_hd__nor2_1 _06349_ (.A(_00490_),
    .B(_00484_),
    .Y(_00491_));
 sky130_fd_sc_hd__nand2_1 _06350_ (.A(_00484_),
    .B(_00490_),
    .Y(_00492_));
 sky130_fd_sc_hd__or2b_1 _06351_ (.A(_00491_),
    .B_N(_00492_),
    .X(_00493_));
 sky130_fd_sc_hd__nand2_1 _06352_ (.A(_06285_),
    .B(_00493_),
    .Y(_00494_));
 sky130_fd_sc_hd__a32o_1 _06353_ (.A1(_00489_),
    .A2(_00475_),
    .A3(_00494_),
    .B1(\next_PC[3] ),
    .B2(_00478_),
    .X(_00017_));
 sky130_fd_sc_hd__nand2_1 _06354_ (.A(_00491_),
    .B(\next_PC[4] ),
    .Y(_00495_));
 sky130_fd_sc_hd__or2_1 _06355_ (.A(\next_PC[4] ),
    .B(_00491_),
    .X(_00496_));
 sky130_fd_sc_hd__a21bo_1 _06356_ (.A1(_00495_),
    .A2(_00496_),
    .B1_N(_00486_),
    .X(_00497_));
 sky130_fd_sc_hd__clkbuf_8 _06357_ (.A(\R1[0] ),
    .X(_00498_));
 sky130_fd_sc_hd__or2_1 _06358_ (.A(_00498_),
    .B(_00486_),
    .X(_00499_));
 sky130_fd_sc_hd__a32o_1 _06359_ (.A1(_00497_),
    .A2(_00475_),
    .A3(_00499_),
    .B1(\next_PC[4] ),
    .B2(_00478_),
    .X(_00018_));
 sky130_fd_sc_hd__inv_2 _06360_ (.A(\next_PC[5] ),
    .Y(_00500_));
 sky130_fd_sc_hd__or2_1 _06361_ (.A(_00500_),
    .B(_00495_),
    .X(_00501_));
 sky130_fd_sc_hd__nand2_1 _06362_ (.A(_00495_),
    .B(_00500_),
    .Y(_00502_));
 sky130_fd_sc_hd__a21bo_1 _06363_ (.A1(_00501_),
    .A2(_00502_),
    .B1_N(_00486_),
    .X(_00503_));
 sky130_fd_sc_hd__or2_1 _06364_ (.A(\R1[1] ),
    .B(_00486_),
    .X(_00504_));
 sky130_fd_sc_hd__a32o_1 _06365_ (.A1(_00503_),
    .A2(_00475_),
    .A3(_00504_),
    .B1(\next_PC[5] ),
    .B2(_00478_),
    .X(_00019_));
 sky130_fd_sc_hd__or2_1 _06366_ (.A(\im_reg[6] ),
    .B(_06285_),
    .X(_00505_));
 sky130_fd_sc_hd__inv_2 _06367_ (.A(\next_PC[6] ),
    .Y(_00506_));
 sky130_fd_sc_hd__or2_1 _06368_ (.A(_00506_),
    .B(_00501_),
    .X(_00507_));
 sky130_fd_sc_hd__inv_2 _06369_ (.A(_00507_),
    .Y(_00508_));
 sky130_fd_sc_hd__and2_1 _06370_ (.A(_00501_),
    .B(_00506_),
    .X(_00509_));
 sky130_fd_sc_hd__o21ai_1 _06371_ (.A1(_00508_),
    .A2(_00509_),
    .B1(_06285_),
    .Y(_00510_));
 sky130_fd_sc_hd__a32o_1 _06372_ (.A1(_00505_),
    .A2(_00475_),
    .A3(_00510_),
    .B1(\next_PC[6] ),
    .B2(_00478_),
    .X(_00020_));
 sky130_fd_sc_hd__nand2_1 _06373_ (.A(_00508_),
    .B(\next_PC[7] ),
    .Y(_00511_));
 sky130_fd_sc_hd__or2_1 _06374_ (.A(\next_PC[7] ),
    .B(_00508_),
    .X(_00512_));
 sky130_fd_sc_hd__a21bo_1 _06375_ (.A1(_00511_),
    .A2(_00512_),
    .B1_N(_00486_),
    .X(_00513_));
 sky130_fd_sc_hd__or2_1 _06376_ (.A(\im_reg[7] ),
    .B(_00486_),
    .X(_00514_));
 sky130_fd_sc_hd__a32o_1 _06377_ (.A1(_00513_),
    .A2(_00475_),
    .A3(_00514_),
    .B1(\next_PC[7] ),
    .B2(_00478_),
    .X(_00021_));
 sky130_fd_sc_hd__inv_2 _06378_ (.A(\next_PC[8] ),
    .Y(_00515_));
 sky130_fd_sc_hd__or2_1 _06379_ (.A(_00515_),
    .B(_00511_),
    .X(_00516_));
 sky130_fd_sc_hd__nand2_1 _06380_ (.A(_00511_),
    .B(_00515_),
    .Y(_00517_));
 sky130_fd_sc_hd__a21bo_1 _06381_ (.A1(_00516_),
    .A2(_00517_),
    .B1_N(_00486_),
    .X(_00518_));
 sky130_fd_sc_hd__or2_1 _06382_ (.A(\im_reg[8] ),
    .B(_00486_),
    .X(_00519_));
 sky130_fd_sc_hd__a32o_1 _06383_ (.A1(_00518_),
    .A2(_00475_),
    .A3(_00519_),
    .B1(\next_PC[8] ),
    .B2(_00478_),
    .X(_00022_));
 sky130_fd_sc_hd__or2_1 _06384_ (.A(\im_reg[9] ),
    .B(_06285_),
    .X(_00520_));
 sky130_fd_sc_hd__xor2_1 _06385_ (.A(\next_PC[9] ),
    .B(_00516_),
    .X(_00521_));
 sky130_fd_sc_hd__nand2_1 _06386_ (.A(_06285_),
    .B(_00521_),
    .Y(_00522_));
 sky130_fd_sc_hd__a32o_1 _06387_ (.A1(_00520_),
    .A2(_00475_),
    .A3(_00522_),
    .B1(\next_PC[9] ),
    .B2(_00478_),
    .X(_00023_));
 sky130_fd_sc_hd__inv_2 _06388_ (.A(Qreg2),
    .Y(_00523_));
 sky130_fd_sc_hd__nor2_4 _06389_ (.A(Oreg2),
    .B(Hreg2),
    .Y(_00524_));
 sky130_fd_sc_hd__clkinv_4 _06390_ (.A(_00524_),
    .Y(_00525_));
 sky130_fd_sc_hd__nor2_2 _06391_ (.A(_00523_),
    .B(_00525_),
    .Y(_00526_));
 sky130_fd_sc_hd__inv_2 _06392_ (.A(_00526_),
    .Y(_00527_));
 sky130_fd_sc_hd__inv_2 _06393_ (.A(CMD_multiplication),
    .Y(_00528_));
 sky130_fd_sc_hd__inv_2 _06394_ (.A(_00471_),
    .Y(_00529_));
 sky130_fd_sc_hd__nor2_2 _06395_ (.A(\current_state[5] ),
    .B(_00529_),
    .Y(_00530_));
 sky130_fd_sc_hd__inv_2 _06396_ (.A(_00530_),
    .Y(_00531_));
 sky130_fd_sc_hd__nor2_2 _06397_ (.A(_00528_),
    .B(_00531_),
    .Y(_00532_));
 sky130_fd_sc_hd__inv_2 _06398_ (.A(_00532_),
    .Y(_00533_));
 sky130_fd_sc_hd__nor2_4 _06399_ (.A(_00527_),
    .B(_00533_),
    .Y(_00534_));
 sky130_fd_sc_hd__clkbuf_4 _06400_ (.A(_00534_),
    .X(_00535_));
 sky130_fd_sc_hd__inv_2 _06401_ (.A(\Add.sub ),
    .Y(_00536_));
 sky130_fd_sc_hd__or4_4 _06402_ (.A(_00536_),
    .B(CMD_addition),
    .C(_06264_),
    .D(_00529_),
    .X(_00537_));
 sky130_fd_sc_hd__inv_2 _06403_ (.A(_00537_),
    .Y(_00538_));
 sky130_fd_sc_hd__nand2_1 _06404_ (.A(_00538_),
    .B(_00526_),
    .Y(_00539_));
 sky130_fd_sc_hd__buf_2 _06405_ (.A(_00539_),
    .X(_00540_));
 sky130_fd_sc_hd__clkbuf_4 _06406_ (.A(_00540_),
    .X(_00541_));
 sky130_fd_sc_hd__inv_2 _06407_ (.A(\result_reg_add[0] ),
    .Y(_00542_));
 sky130_fd_sc_hd__a21oi_1 _06408_ (.A1(_00541_),
    .A2(_00542_),
    .B1(_00535_),
    .Y(_00543_));
 sky130_fd_sc_hd__or2_1 _06409_ (.A(\result_reg_sub[0] ),
    .B(_00540_),
    .X(_00544_));
 sky130_fd_sc_hd__clkbuf_4 _06410_ (.A(CMD_or),
    .X(_00545_));
 sky130_fd_sc_hd__nor2_1 _06411_ (.A(\shift.left ),
    .B(CMD_logic_shift_right),
    .Y(_00546_));
 sky130_fd_sc_hd__inv_2 _06412_ (.A(CMD_and),
    .Y(_00547_));
 sky130_fd_sc_hd__inv_2 _06413_ (.A(CMD_mul_accumulation),
    .Y(_00548_));
 sky130_fd_sc_hd__buf_4 _06414_ (.A(_00548_),
    .X(_00549_));
 sky130_fd_sc_hd__and3_2 _06415_ (.A(_00546_),
    .B(_00547_),
    .C(_00549_),
    .X(_00550_));
 sky130_fd_sc_hd__and4_2 _06416_ (.A(_00530_),
    .B(_00545_),
    .C(_00528_),
    .D(_00550_),
    .X(_00551_));
 sky130_fd_sc_hd__nand2_2 _06417_ (.A(_00551_),
    .B(_00526_),
    .Y(_00552_));
 sky130_fd_sc_hd__buf_2 _06418_ (.A(_00552_),
    .X(_00553_));
 sky130_fd_sc_hd__inv_2 _06419_ (.A(_00546_),
    .Y(_00554_));
 sky130_fd_sc_hd__nor2_1 _06420_ (.A(_00547_),
    .B(_00554_),
    .Y(_00555_));
 sky130_fd_sc_hd__buf_4 _06421_ (.A(_00549_),
    .X(_00556_));
 sky130_fd_sc_hd__clkbuf_4 _06422_ (.A(CMD_multiplication),
    .X(_00557_));
 sky130_fd_sc_hd__nor2_1 _06423_ (.A(_00557_),
    .B(\current_state[5] ),
    .Y(_00558_));
 sky130_fd_sc_hd__and4_2 _06424_ (.A(_00472_),
    .B(_00555_),
    .C(_00556_),
    .D(_00558_),
    .X(_00559_));
 sky130_fd_sc_hd__nand2_1 _06425_ (.A(_00559_),
    .B(_00526_),
    .Y(_00560_));
 sky130_fd_sc_hd__clkbuf_4 _06426_ (.A(_00560_),
    .X(_00561_));
 sky130_fd_sc_hd__clkbuf_4 _06427_ (.A(_00561_),
    .X(_00562_));
 sky130_fd_sc_hd__nand2_1 _06428_ (.A(_00553_),
    .B(_00562_),
    .Y(_00563_));
 sky130_fd_sc_hd__a221o_1 _06429_ (.A1(\result_reg_mul[0] ),
    .A2(_00535_),
    .B1(_00543_),
    .B2(_00544_),
    .C1(_00563_),
    .X(_00564_));
 sky130_fd_sc_hd__and3_1 _06430_ (.A(_00471_),
    .B(CMD_addition),
    .C(\current_state[5] ),
    .X(_00565_));
 sky130_fd_sc_hd__inv_2 _06431_ (.A(_00565_),
    .Y(_00566_));
 sky130_fd_sc_hd__nand2_1 _06432_ (.A(_00533_),
    .B(_00566_),
    .Y(_00567_));
 sky130_fd_sc_hd__nor2_2 _06433_ (.A(_00567_),
    .B(_00538_),
    .Y(_00568_));
 sky130_fd_sc_hd__inv_2 _06434_ (.A(_00568_),
    .Y(_00569_));
 sky130_fd_sc_hd__inv_2 _06435_ (.A(Oim),
    .Y(_00570_));
 sky130_fd_sc_hd__nand2_1 _06436_ (.A(_00570_),
    .B(Qim),
    .Y(_00571_));
 sky130_fd_sc_hd__nor2_2 _06437_ (.A(Qreg2),
    .B(_00525_),
    .Y(_00572_));
 sky130_fd_sc_hd__inv_2 _06438_ (.A(_00572_),
    .Y(_00573_));
 sky130_fd_sc_hd__nor3_4 _06439_ (.A(Him),
    .B(_00571_),
    .C(_00573_),
    .Y(_00574_));
 sky130_fd_sc_hd__nand2_1 _06440_ (.A(_00569_),
    .B(_00574_),
    .Y(_00575_));
 sky130_fd_sc_hd__inv_2 _06441_ (.A(CMD_set),
    .Y(_00576_));
 sky130_fd_sc_hd__nor2_1 _06442_ (.A(_00545_),
    .B(_00576_),
    .Y(_00577_));
 sky130_fd_sc_hd__inv_2 _06443_ (.A(CMD_not),
    .Y(_00578_));
 sky130_fd_sc_hd__nand2_1 _06444_ (.A(_00577_),
    .B(_00578_),
    .Y(_00579_));
 sky130_fd_sc_hd__inv_2 _06445_ (.A(\shift.Q ),
    .Y(_00580_));
 sky130_fd_sc_hd__clkbuf_4 _06446_ (.A(_00580_),
    .X(_00581_));
 sky130_fd_sc_hd__buf_4 _06447_ (.A(_00581_),
    .X(_00582_));
 sky130_fd_sc_hd__buf_4 _06448_ (.A(\shift.O ),
    .X(_00583_));
 sky130_fd_sc_hd__clkbuf_4 _06449_ (.A(_00583_),
    .X(_00584_));
 sky130_fd_sc_hd__buf_4 _06450_ (.A(_00584_),
    .X(_00585_));
 sky130_fd_sc_hd__buf_6 _06451_ (.A(\shift.H ),
    .X(_00586_));
 sky130_fd_sc_hd__buf_6 _06452_ (.A(_00586_),
    .X(_00587_));
 sky130_fd_sc_hd__clkbuf_4 _06453_ (.A(_00587_),
    .X(_00588_));
 sky130_fd_sc_hd__buf_4 _06454_ (.A(_00588_),
    .X(_00589_));
 sky130_fd_sc_hd__nor2_4 _06455_ (.A(_00585_),
    .B(_00589_),
    .Y(_00590_));
 sky130_fd_sc_hd__inv_4 _06456_ (.A(_00590_),
    .Y(_00591_));
 sky130_fd_sc_hd__nor2_2 _06457_ (.A(_00582_),
    .B(_00591_),
    .Y(_00592_));
 sky130_fd_sc_hd__inv_2 _06458_ (.A(_00592_),
    .Y(_00593_));
 sky130_fd_sc_hd__nor2_1 _06459_ (.A(_00593_),
    .B(_00531_),
    .Y(_00594_));
 sky130_fd_sc_hd__and3_1 _06460_ (.A(_00594_),
    .B(_00528_),
    .C(_00550_),
    .X(_00595_));
 sky130_fd_sc_hd__or2b_1 _06461_ (.A(_00579_),
    .B_N(_00595_),
    .X(_00596_));
 sky130_fd_sc_hd__nor2_1 _06462_ (.A(CMD_set),
    .B(_00545_),
    .Y(_00597_));
 sky130_fd_sc_hd__and3_1 _06463_ (.A(_00597_),
    .B(CMD_load),
    .C(_00578_),
    .X(_00598_));
 sky130_fd_sc_hd__and2_1 _06464_ (.A(_00595_),
    .B(_00598_),
    .X(_00599_));
 sky130_fd_sc_hd__buf_2 _06465_ (.A(_00599_),
    .X(_00600_));
 sky130_fd_sc_hd__inv_2 _06466_ (.A(_00600_),
    .Y(_00601_));
 sky130_fd_sc_hd__and3_1 _06467_ (.A(_00575_),
    .B(_00596_),
    .C(_00601_),
    .X(_00602_));
 sky130_fd_sc_hd__clkbuf_4 _06468_ (.A(_00602_),
    .X(_00603_));
 sky130_fd_sc_hd__o221a_1 _06469_ (.A1(\result_reg_or[0] ),
    .A2(_00553_),
    .B1(\result_reg_and[0] ),
    .B2(_00562_),
    .C1(_00603_),
    .X(_00604_));
 sky130_fd_sc_hd__nand2_1 _06470_ (.A(_00550_),
    .B(_00592_),
    .Y(_00605_));
 sky130_fd_sc_hd__nand2_1 _06471_ (.A(_00530_),
    .B(_00528_),
    .Y(_00606_));
 sky130_fd_sc_hd__or3_2 _06472_ (.A(_00579_),
    .B(_00605_),
    .C(_00606_),
    .X(_00607_));
 sky130_fd_sc_hd__clkbuf_4 _06473_ (.A(_00607_),
    .X(_00608_));
 sky130_fd_sc_hd__inv_2 _06474_ (.A(\result_reg_mul[0] ),
    .Y(_00609_));
 sky130_fd_sc_hd__inv_2 _06475_ (.A(\result_reg_sub[0] ),
    .Y(_00610_));
 sky130_fd_sc_hd__nand2_4 _06476_ (.A(_00538_),
    .B(_00574_),
    .Y(_00611_));
 sky130_fd_sc_hd__mux2_1 _06477_ (.A0(_00610_),
    .A1(_00542_),
    .S(_00611_),
    .X(_00612_));
 sky130_fd_sc_hd__nand2_4 _06478_ (.A(_00532_),
    .B(_00574_),
    .Y(_00613_));
 sky130_fd_sc_hd__mux2_1 _06479_ (.A0(_00609_),
    .A1(_00612_),
    .S(_00613_),
    .X(_00614_));
 sky130_fd_sc_hd__buf_2 _06480_ (.A(_00607_),
    .X(_00615_));
 sky130_fd_sc_hd__nand2_1 _06481_ (.A(_00614_),
    .B(_00615_),
    .Y(_00616_));
 sky130_fd_sc_hd__o211a_1 _06482_ (.A1(\result_reg_set[0] ),
    .A2(_00608_),
    .B1(_00601_),
    .C1(_00616_),
    .X(_00617_));
 sky130_fd_sc_hd__a21o_1 _06483_ (.A1(net1),
    .A2(_00600_),
    .B1(_00617_),
    .X(_00618_));
 sky130_fd_sc_hd__inv_2 _06484_ (.A(_00603_),
    .Y(_00619_));
 sky130_fd_sc_hd__inv_2 _06485_ (.A(Qreg3),
    .Y(_00620_));
 sky130_fd_sc_hd__clkbuf_8 _06486_ (.A(Oreg3),
    .X(_00621_));
 sky130_fd_sc_hd__clkbuf_4 _06487_ (.A(CMD_mul_accumulation),
    .X(_00622_));
 sky130_fd_sc_hd__clkbuf_4 _06488_ (.A(_00622_),
    .X(_00623_));
 sky130_fd_sc_hd__buf_4 _06489_ (.A(_00623_),
    .X(_00624_));
 sky130_fd_sc_hd__nand2_2 _06490_ (.A(_00558_),
    .B(_00624_),
    .Y(_00625_));
 sky130_fd_sc_hd__inv_4 _06491_ (.A(Hreg3),
    .Y(_00626_));
 sky130_fd_sc_hd__nand2_1 _06492_ (.A(_00472_),
    .B(_00626_),
    .Y(_00627_));
 sky130_fd_sc_hd__or4_4 _06493_ (.A(_00620_),
    .B(_00621_),
    .C(_00625_),
    .D(_00627_),
    .X(_00628_));
 sky130_fd_sc_hd__inv_2 _06494_ (.A(_00628_),
    .Y(_00629_));
 sky130_fd_sc_hd__a221o_1 _06495_ (.A1(_00564_),
    .A2(_00604_),
    .B1(_00618_),
    .B2(_00619_),
    .C1(_00629_),
    .X(_00630_));
 sky130_fd_sc_hd__buf_2 _06496_ (.A(\current_state[5] ),
    .X(_00631_));
 sky130_fd_sc_hd__or3_4 _06497_ (.A(CMD_or),
    .B(CMD_multiplication),
    .C(_00578_),
    .X(_00632_));
 sky130_fd_sc_hd__nor2_2 _06498_ (.A(_00631_),
    .B(_00632_),
    .Y(_00633_));
 sky130_fd_sc_hd__buf_2 _06499_ (.A(_00529_),
    .X(_00634_));
 sky130_fd_sc_hd__buf_4 _06500_ (.A(_00634_),
    .X(_00635_));
 sky130_fd_sc_hd__nor2_2 _06501_ (.A(_00635_),
    .B(_00605_),
    .Y(_00636_));
 sky130_fd_sc_hd__inv_2 _06502_ (.A(CMD_logic_shift_right),
    .Y(_00637_));
 sky130_fd_sc_hd__nor2_1 _06503_ (.A(_00623_),
    .B(_00557_),
    .Y(_00638_));
 sky130_fd_sc_hd__inv_2 _06504_ (.A(_00638_),
    .Y(_00639_));
 sky130_fd_sc_hd__nor2_2 _06505_ (.A(_00637_),
    .B(_00639_),
    .Y(_00640_));
 sky130_fd_sc_hd__and3_2 _06506_ (.A(_00638_),
    .B(\shift.left ),
    .C(_00637_),
    .X(_00641_));
 sky130_fd_sc_hd__and3_1 _06507_ (.A(_00530_),
    .B(_00592_),
    .C(_00641_),
    .X(_00642_));
 sky130_fd_sc_hd__buf_4 _06508_ (.A(_00642_),
    .X(_00643_));
 sky130_fd_sc_hd__a221o_4 _06509_ (.A1(_00633_),
    .A2(_00636_),
    .B1(_00594_),
    .B2(_00640_),
    .C1(_00643_),
    .X(_00644_));
 sky130_fd_sc_hd__inv_2 _06510_ (.A(_00644_),
    .Y(_00645_));
 sky130_fd_sc_hd__inv_2 _06511_ (.A(Oreg3),
    .Y(_00646_));
 sky130_fd_sc_hd__clkbuf_8 _06512_ (.A(_00646_),
    .X(_00647_));
 sky130_fd_sc_hd__and3_1 _06513_ (.A(_00647_),
    .B(_00626_),
    .C(Qreg3),
    .X(_00648_));
 sky130_fd_sc_hd__and3b_1 _06514_ (.A_N(_00625_),
    .B(_00472_),
    .C(_00648_),
    .X(_00649_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06515_ (.A(_00649_),
    .X(_00650_));
 sky130_fd_sc_hd__or2b_1 _06516_ (.A(\result_reg_mac[0] ),
    .B_N(_00650_),
    .X(_00651_));
 sky130_fd_sc_hd__inv_2 _06517_ (.A(\result_reg_not[0] ),
    .Y(_00652_));
 sky130_fd_sc_hd__inv_2 _06518_ (.A(_00550_),
    .Y(_00653_));
 sky130_fd_sc_hd__nor2_8 _06519_ (.A(_00632_),
    .B(_00653_),
    .Y(_00654_));
 sky130_fd_sc_hd__clkbuf_4 _06520_ (.A(_00654_),
    .X(_00655_));
 sky130_fd_sc_hd__nand2_4 _06521_ (.A(_00636_),
    .B(_00633_),
    .Y(_00656_));
 sky130_fd_sc_hd__clkbuf_4 _06522_ (.A(_00656_),
    .X(_00657_));
 sky130_fd_sc_hd__inv_2 _06523_ (.A(\result_reg_Rshift[0] ),
    .Y(_00658_));
 sky130_fd_sc_hd__inv_2 _06524_ (.A(\result_reg_Lshift[0] ),
    .Y(_00659_));
 sky130_fd_sc_hd__mux2_1 _06525_ (.A0(_00658_),
    .A1(_00659_),
    .S(_00643_),
    .X(_00660_));
 sky130_fd_sc_hd__nor2_2 _06526_ (.A(_00546_),
    .B(_00639_),
    .Y(_00661_));
 sky130_fd_sc_hd__inv_2 _06527_ (.A(_00545_),
    .Y(_00662_));
 sky130_fd_sc_hd__and3_1 _06528_ (.A(_00595_),
    .B(CMD_not),
    .C(_00662_),
    .X(_00663_));
 sky130_fd_sc_hd__a21o_4 _06529_ (.A1(_00594_),
    .A2(_00661_),
    .B1(_00663_),
    .X(_00664_));
 sky130_fd_sc_hd__clkinv_4 _06530_ (.A(_00664_),
    .Y(_00665_));
 sky130_fd_sc_hd__clkbuf_4 _06531_ (.A(_00665_),
    .X(_00666_));
 sky130_fd_sc_hd__a221oi_2 _06532_ (.A1(_00652_),
    .A2(_00655_),
    .B1(_00657_),
    .B2(_00660_),
    .C1(_00666_),
    .Y(_00667_));
 sky130_fd_sc_hd__a31o_2 _06533_ (.A1(_00630_),
    .A2(_00645_),
    .A3(_00651_),
    .B1(_00667_),
    .X(_00668_));
 sky130_fd_sc_hd__inv_2 _06534_ (.A(\R3[1] ),
    .Y(_00669_));
 sky130_fd_sc_hd__inv_2 _06535_ (.A(\R0[1] ),
    .Y(_00670_));
 sky130_fd_sc_hd__inv_2 _06536_ (.A(\R2[1] ),
    .Y(_00671_));
 sky130_fd_sc_hd__mux2_1 _06537_ (.A0(_00670_),
    .A1(_00671_),
    .S(_00602_),
    .X(_00672_));
 sky130_fd_sc_hd__nor2_1 _06538_ (.A(\R1[1] ),
    .B(_00628_),
    .Y(_00673_));
 sky130_fd_sc_hd__a211o_1 _06539_ (.A1(_00672_),
    .A2(_00628_),
    .B1(_00664_),
    .C1(_00673_),
    .X(_00674_));
 sky130_fd_sc_hd__o21a_1 _06540_ (.A1(_00669_),
    .A2(_00665_),
    .B1(_00674_),
    .X(_00675_));
 sky130_fd_sc_hd__and3_1 _06541_ (.A(_00628_),
    .B(_00560_),
    .C(_00552_),
    .X(_00676_));
 sky130_fd_sc_hd__o2111ai_4 _06542_ (.A1(_00568_),
    .A2(_00527_),
    .B1(_00665_),
    .C1(_00676_),
    .D1(_00603_),
    .Y(_00677_));
 sky130_fd_sc_hd__nand2_1 _06543_ (.A(_00675_),
    .B(_00677_),
    .Y(_00678_));
 sky130_fd_sc_hd__inv_2 _06544_ (.A(_00678_),
    .Y(_00679_));
 sky130_fd_sc_hd__o21a_1 _06545_ (.A1(\R0[0] ),
    .A2(_00602_),
    .B1(_00628_),
    .X(_00680_));
 sky130_fd_sc_hd__inv_2 _06546_ (.A(\R2[0] ),
    .Y(_00681_));
 sky130_fd_sc_hd__nand2_1 _06547_ (.A(_00602_),
    .B(_00681_),
    .Y(_00682_));
 sky130_fd_sc_hd__a221o_1 _06548_ (.A1(_00498_),
    .A2(_00629_),
    .B1(_00680_),
    .B2(_00682_),
    .C1(_00664_),
    .X(_00683_));
 sky130_fd_sc_hd__o21a_1 _06549_ (.A1(\R3[0] ),
    .A2(_00665_),
    .B1(_00683_),
    .X(_00684_));
 sky130_fd_sc_hd__inv_2 _06550_ (.A(_00684_),
    .Y(_00685_));
 sky130_fd_sc_hd__nand2_4 _06551_ (.A(_00679_),
    .B(_00685_),
    .Y(_00686_));
 sky130_fd_sc_hd__buf_6 _06552_ (.A(_00686_),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _06553_ (.A0(_00668_),
    .A1(\Qset[0][0] ),
    .S(_00687_),
    .X(_00688_));
 sky130_fd_sc_hd__clkbuf_1 _06554_ (.A(_00688_),
    .X(_00024_));
 sky130_fd_sc_hd__inv_2 _06555_ (.A(\result_reg_not[1] ),
    .Y(_00689_));
 sky130_fd_sc_hd__inv_2 _06556_ (.A(\result_reg_Rshift[1] ),
    .Y(_00690_));
 sky130_fd_sc_hd__inv_2 _06557_ (.A(\result_reg_Lshift[1] ),
    .Y(_00691_));
 sky130_fd_sc_hd__mux2_1 _06558_ (.A0(_00690_),
    .A1(_00691_),
    .S(_00643_),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _06559_ (.A0(_00689_),
    .A1(_00692_),
    .S(_00656_),
    .X(_00693_));
 sky130_fd_sc_hd__inv_2 _06560_ (.A(\result_reg_mac[1] ),
    .Y(_00694_));
 sky130_fd_sc_hd__clkbuf_4 _06561_ (.A(_00650_),
    .X(_00695_));
 sky130_fd_sc_hd__buf_2 _06562_ (.A(_00601_),
    .X(_00696_));
 sky130_fd_sc_hd__inv_2 _06563_ (.A(CMD_load),
    .Y(_00697_));
 sky130_fd_sc_hd__nand2_1 _06564_ (.A(_00597_),
    .B(_00578_),
    .Y(_00698_));
 sky130_fd_sc_hd__or4_4 _06565_ (.A(_00697_),
    .B(_00605_),
    .C(_00698_),
    .D(_00606_),
    .X(_00699_));
 sky130_fd_sc_hd__inv_2 _06566_ (.A(\result_reg_set[1] ),
    .Y(_00700_));
 sky130_fd_sc_hd__inv_2 _06567_ (.A(\result_reg_mul[1] ),
    .Y(_00701_));
 sky130_fd_sc_hd__inv_2 _06568_ (.A(\result_reg_sub[1] ),
    .Y(_00702_));
 sky130_fd_sc_hd__inv_2 _06569_ (.A(\result_reg_add[1] ),
    .Y(_00703_));
 sky130_fd_sc_hd__mux2_1 _06570_ (.A0(_00702_),
    .A1(_00703_),
    .S(_00611_),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _06571_ (.A0(_00701_),
    .A1(_00704_),
    .S(_00613_),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_1 _06572_ (.A0(_00700_),
    .A1(_00705_),
    .S(_00607_),
    .X(_00706_));
 sky130_fd_sc_hd__a2bb2o_1 _06573_ (.A1_N(net8),
    .A2_N(_00696_),
    .B1(_00699_),
    .B2(_00706_),
    .X(_00707_));
 sky130_fd_sc_hd__inv_2 _06574_ (.A(\result_reg_or[1] ),
    .Y(_00708_));
 sky130_fd_sc_hd__buf_2 _06575_ (.A(_00552_),
    .X(_00709_));
 sky130_fd_sc_hd__buf_6 _06576_ (.A(_00624_),
    .X(_00710_));
 sky130_fd_sc_hd__or3_1 _06577_ (.A(_00662_),
    .B(CMD_and),
    .C(_00527_),
    .X(_00711_));
 sky130_fd_sc_hd__or4_1 _06578_ (.A(\shift.left ),
    .B(CMD_logic_shift_right),
    .C(_00710_),
    .D(_00711_),
    .X(_00712_));
 sky130_fd_sc_hd__or4_1 _06579_ (.A(_00557_),
    .B(_00631_),
    .C(_00634_),
    .D(_00712_),
    .X(_00713_));
 sky130_fd_sc_hd__inv_2 _06580_ (.A(_00713_),
    .Y(_00714_));
 sky130_fd_sc_hd__inv_2 _06581_ (.A(\result_reg_and[1] ),
    .Y(_00715_));
 sky130_fd_sc_hd__mux2_1 _06582_ (.A0(_00702_),
    .A1(_00703_),
    .S(_00539_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _06583_ (.A0(_00716_),
    .A1(_00701_),
    .S(_00534_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _06584_ (.A0(_00715_),
    .A1(_00717_),
    .S(_00560_),
    .X(_00718_));
 sky130_fd_sc_hd__o221a_1 _06585_ (.A1(_00708_),
    .A2(_00709_),
    .B1(_00714_),
    .B2(_00718_),
    .C1(_00603_),
    .X(_00719_));
 sky130_fd_sc_hd__a21o_1 _06586_ (.A1(_00707_),
    .A2(_00619_),
    .B1(_00719_),
    .X(_00720_));
 sky130_fd_sc_hd__a221o_1 _06587_ (.A1(_00694_),
    .A2(_00695_),
    .B1(_00720_),
    .B2(_00628_),
    .C1(_00644_),
    .X(_00721_));
 sky130_fd_sc_hd__o21ai_4 _06588_ (.A1(_00645_),
    .A2(_00693_),
    .B1(_00721_),
    .Y(_00722_));
 sky130_fd_sc_hd__mux2_1 _06589_ (.A0(_00722_),
    .A1(\Qset[0][1] ),
    .S(_00687_),
    .X(_00723_));
 sky130_fd_sc_hd__clkbuf_1 _06590_ (.A(_00723_),
    .X(_00025_));
 sky130_fd_sc_hd__inv_2 _06591_ (.A(\result_reg_mac[2] ),
    .Y(_00724_));
 sky130_fd_sc_hd__clkbuf_4 _06592_ (.A(_00628_),
    .X(_00725_));
 sky130_fd_sc_hd__inv_2 _06593_ (.A(\result_reg_set[2] ),
    .Y(_00726_));
 sky130_fd_sc_hd__inv_2 _06594_ (.A(\result_reg_mul[2] ),
    .Y(_00727_));
 sky130_fd_sc_hd__inv_2 _06595_ (.A(\result_reg_sub[2] ),
    .Y(_00728_));
 sky130_fd_sc_hd__inv_2 _06596_ (.A(\result_reg_add[2] ),
    .Y(_00729_));
 sky130_fd_sc_hd__buf_4 _06597_ (.A(_00611_),
    .X(_00730_));
 sky130_fd_sc_hd__mux2_1 _06598_ (.A0(_00728_),
    .A1(_00729_),
    .S(_00730_),
    .X(_00731_));
 sky130_fd_sc_hd__clkbuf_4 _06599_ (.A(_00613_),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_1 _06600_ (.A0(_00727_),
    .A1(_00731_),
    .S(_00732_),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _06601_ (.A0(_00726_),
    .A1(_00733_),
    .S(_00608_),
    .X(_00734_));
 sky130_fd_sc_hd__clkbuf_4 _06602_ (.A(_00699_),
    .X(_00735_));
 sky130_fd_sc_hd__nand2_1 _06603_ (.A(_00734_),
    .B(_00735_),
    .Y(_00736_));
 sky130_fd_sc_hd__o21ai_1 _06604_ (.A1(net9),
    .A2(_00696_),
    .B1(_00736_),
    .Y(_00737_));
 sky130_fd_sc_hd__inv_2 _06605_ (.A(\result_reg_or[2] ),
    .Y(_00738_));
 sky130_fd_sc_hd__buf_2 _06606_ (.A(_00603_),
    .X(_00739_));
 sky130_fd_sc_hd__clkbuf_4 _06607_ (.A(_00540_),
    .X(_00740_));
 sky130_fd_sc_hd__a21oi_1 _06608_ (.A1(_00540_),
    .A2(_00729_),
    .B1(_00534_),
    .Y(_00741_));
 sky130_fd_sc_hd__o21ai_1 _06609_ (.A1(\result_reg_sub[2] ),
    .A2(_00740_),
    .B1(_00741_),
    .Y(_00742_));
 sky130_fd_sc_hd__buf_2 _06610_ (.A(_00561_),
    .X(_00743_));
 sky130_fd_sc_hd__or4_2 _06611_ (.A(_00528_),
    .B(_00631_),
    .C(_00527_),
    .D(_00634_),
    .X(_00744_));
 sky130_fd_sc_hd__clkbuf_2 _06612_ (.A(_00744_),
    .X(_00745_));
 sky130_fd_sc_hd__or2_1 _06613_ (.A(_00727_),
    .B(_00745_),
    .X(_00746_));
 sky130_fd_sc_hd__o21ai_2 _06614_ (.A1(\result_reg_and[2] ),
    .A2(_00561_),
    .B1(_00552_),
    .Y(_00747_));
 sky130_fd_sc_hd__a31o_1 _06615_ (.A1(_00742_),
    .A2(_00743_),
    .A3(_00746_),
    .B1(_00747_),
    .X(_00748_));
 sky130_fd_sc_hd__o211a_1 _06616_ (.A1(_00738_),
    .A2(_00709_),
    .B1(_00739_),
    .C1(_00748_),
    .X(_00749_));
 sky130_fd_sc_hd__a211o_1 _06617_ (.A1(_00737_),
    .A2(_00619_),
    .B1(_00629_),
    .C1(_00749_),
    .X(_00750_));
 sky130_fd_sc_hd__o21a_1 _06618_ (.A1(_00724_),
    .A2(_00725_),
    .B1(_00750_),
    .X(_00751_));
 sky130_fd_sc_hd__inv_2 _06619_ (.A(\result_reg_not[2] ),
    .Y(_00752_));
 sky130_fd_sc_hd__clkbuf_4 _06620_ (.A(_00643_),
    .X(_00753_));
 sky130_fd_sc_hd__buf_2 _06621_ (.A(_00643_),
    .X(_00754_));
 sky130_fd_sc_hd__inv_2 _06622_ (.A(\result_reg_Lshift[2] ),
    .Y(_00755_));
 sky130_fd_sc_hd__nand2_1 _06623_ (.A(_00754_),
    .B(_00755_),
    .Y(_00756_));
 sky130_fd_sc_hd__o21ai_1 _06624_ (.A1(\result_reg_Rshift[2] ),
    .A2(_00753_),
    .B1(_00756_),
    .Y(_00757_));
 sky130_fd_sc_hd__a221o_2 _06625_ (.A1(_00752_),
    .A2(_00655_),
    .B1(_00657_),
    .B2(_00757_),
    .C1(_00666_),
    .X(_00758_));
 sky130_fd_sc_hd__o21ai_4 _06626_ (.A1(_00664_),
    .A2(_00751_),
    .B1(_00758_),
    .Y(_00759_));
 sky130_fd_sc_hd__mux2_1 _06627_ (.A0(_00759_),
    .A1(\Qset[0][2] ),
    .S(_00687_),
    .X(_00760_));
 sky130_fd_sc_hd__clkbuf_1 _06628_ (.A(_00760_),
    .X(_00026_));
 sky130_fd_sc_hd__inv_2 _06629_ (.A(\result_reg_mac[3] ),
    .Y(_00761_));
 sky130_fd_sc_hd__inv_2 _06630_ (.A(\result_reg_add[3] ),
    .Y(_00762_));
 sky130_fd_sc_hd__a21oi_1 _06631_ (.A1(_00740_),
    .A2(_00762_),
    .B1(_00535_),
    .Y(_00763_));
 sky130_fd_sc_hd__o21ai_1 _06632_ (.A1(\result_reg_sub[3] ),
    .A2(_00541_),
    .B1(_00763_),
    .Y(_00764_));
 sky130_fd_sc_hd__inv_2 _06633_ (.A(\result_reg_mul[3] ),
    .Y(_00765_));
 sky130_fd_sc_hd__or2_1 _06634_ (.A(_00765_),
    .B(_00745_),
    .X(_00766_));
 sky130_fd_sc_hd__o21ai_1 _06635_ (.A1(\result_reg_and[3] ),
    .A2(_00743_),
    .B1(_00553_),
    .Y(_00767_));
 sky130_fd_sc_hd__a31o_1 _06636_ (.A1(_00764_),
    .A2(_00562_),
    .A3(_00766_),
    .B1(_00767_),
    .X(_00768_));
 sky130_fd_sc_hd__or2b_1 _06637_ (.A(_00553_),
    .B_N(\result_reg_or[3] ),
    .X(_00769_));
 sky130_fd_sc_hd__inv_2 _06638_ (.A(\result_reg_sub[3] ),
    .Y(_00770_));
 sky130_fd_sc_hd__mux2_1 _06639_ (.A0(_00770_),
    .A1(_00762_),
    .S(_00730_),
    .X(_00771_));
 sky130_fd_sc_hd__mux2_1 _06640_ (.A0(_00765_),
    .A1(_00771_),
    .S(_00732_),
    .X(_00772_));
 sky130_fd_sc_hd__nand2_1 _06641_ (.A(_00772_),
    .B(_00615_),
    .Y(_00773_));
 sky130_fd_sc_hd__o211ai_1 _06642_ (.A1(\result_reg_set[3] ),
    .A2(_00615_),
    .B1(_00696_),
    .C1(_00773_),
    .Y(_00774_));
 sky130_fd_sc_hd__a21oi_1 _06643_ (.A1(net10),
    .A2(_00600_),
    .B1(_00739_),
    .Y(_00775_));
 sky130_fd_sc_hd__a32o_1 _06644_ (.A1(_00739_),
    .A2(_00768_),
    .A3(_00769_),
    .B1(_00774_),
    .B2(_00775_),
    .X(_00776_));
 sky130_fd_sc_hd__a221o_1 _06645_ (.A1(_00761_),
    .A2(_00695_),
    .B1(_00776_),
    .B2(_00725_),
    .C1(_00644_),
    .X(_00777_));
 sky130_fd_sc_hd__inv_2 _06646_ (.A(\result_reg_not[3] ),
    .Y(_00778_));
 sky130_fd_sc_hd__inv_2 _06647_ (.A(\result_reg_Lshift[3] ),
    .Y(_00779_));
 sky130_fd_sc_hd__nand2_1 _06648_ (.A(_00754_),
    .B(_00779_),
    .Y(_00780_));
 sky130_fd_sc_hd__o21ai_1 _06649_ (.A1(\result_reg_Rshift[3] ),
    .A2(_00753_),
    .B1(_00780_),
    .Y(_00781_));
 sky130_fd_sc_hd__a221o_1 _06650_ (.A1(_00778_),
    .A2(_00655_),
    .B1(_00657_),
    .B2(_00781_),
    .C1(_00666_),
    .X(_00782_));
 sky130_fd_sc_hd__nand2_4 _06651_ (.A(_00777_),
    .B(_00782_),
    .Y(_00783_));
 sky130_fd_sc_hd__mux2_1 _06652_ (.A0(_00783_),
    .A1(\Qset[0][3] ),
    .S(_00687_),
    .X(_00784_));
 sky130_fd_sc_hd__clkbuf_1 _06653_ (.A(_00784_),
    .X(_00027_));
 sky130_fd_sc_hd__inv_2 _06654_ (.A(\result_reg_mac[4] ),
    .Y(_00785_));
 sky130_fd_sc_hd__inv_2 _06655_ (.A(\result_reg_set[4] ),
    .Y(_00786_));
 sky130_fd_sc_hd__inv_2 _06656_ (.A(\result_reg_mul[4] ),
    .Y(_00787_));
 sky130_fd_sc_hd__inv_2 _06657_ (.A(\result_reg_sub[4] ),
    .Y(_00788_));
 sky130_fd_sc_hd__inv_2 _06658_ (.A(\result_reg_add[4] ),
    .Y(_00789_));
 sky130_fd_sc_hd__mux2_1 _06659_ (.A0(_00788_),
    .A1(_00789_),
    .S(_00730_),
    .X(_00790_));
 sky130_fd_sc_hd__mux2_1 _06660_ (.A0(_00787_),
    .A1(_00790_),
    .S(_00732_),
    .X(_00791_));
 sky130_fd_sc_hd__mux2_1 _06661_ (.A0(_00786_),
    .A1(_00791_),
    .S(_00608_),
    .X(_00792_));
 sky130_fd_sc_hd__nand2_1 _06662_ (.A(_00792_),
    .B(_00735_),
    .Y(_00793_));
 sky130_fd_sc_hd__o21ai_1 _06663_ (.A1(net11),
    .A2(_00696_),
    .B1(_00793_),
    .Y(_00794_));
 sky130_fd_sc_hd__inv_2 _06664_ (.A(\result_reg_or[4] ),
    .Y(_00795_));
 sky130_fd_sc_hd__a21oi_1 _06665_ (.A1(_00540_),
    .A2(_00789_),
    .B1(_00534_),
    .Y(_00796_));
 sky130_fd_sc_hd__o21ai_1 _06666_ (.A1(\result_reg_sub[4] ),
    .A2(_00740_),
    .B1(_00796_),
    .Y(_00797_));
 sky130_fd_sc_hd__or2_1 _06667_ (.A(_00787_),
    .B(_00745_),
    .X(_00798_));
 sky130_fd_sc_hd__o21ai_1 _06668_ (.A1(\result_reg_and[4] ),
    .A2(_00561_),
    .B1(_00552_),
    .Y(_00799_));
 sky130_fd_sc_hd__a31o_1 _06669_ (.A1(_00797_),
    .A2(_00743_),
    .A3(_00798_),
    .B1(_00799_),
    .X(_00800_));
 sky130_fd_sc_hd__o211a_1 _06670_ (.A1(_00795_),
    .A2(_00709_),
    .B1(_00739_),
    .C1(_00800_),
    .X(_00801_));
 sky130_fd_sc_hd__a211o_1 _06671_ (.A1(_00794_),
    .A2(_00619_),
    .B1(_00629_),
    .C1(_00801_),
    .X(_00802_));
 sky130_fd_sc_hd__o21a_1 _06672_ (.A1(_00785_),
    .A2(_00725_),
    .B1(_00802_),
    .X(_00803_));
 sky130_fd_sc_hd__inv_2 _06673_ (.A(\result_reg_not[4] ),
    .Y(_00804_));
 sky130_fd_sc_hd__inv_2 _06674_ (.A(\result_reg_Rshift[4] ),
    .Y(_00805_));
 sky130_fd_sc_hd__inv_2 _06675_ (.A(\result_reg_Lshift[4] ),
    .Y(_00806_));
 sky130_fd_sc_hd__mux2_1 _06676_ (.A0(_00805_),
    .A1(_00806_),
    .S(_00643_),
    .X(_00807_));
 sky130_fd_sc_hd__a221o_1 _06677_ (.A1(_00804_),
    .A2(_00655_),
    .B1(_00657_),
    .B2(_00807_),
    .C1(_00666_),
    .X(_00808_));
 sky130_fd_sc_hd__o21ai_4 _06678_ (.A1(_00664_),
    .A2(_00803_),
    .B1(_00808_),
    .Y(_00809_));
 sky130_fd_sc_hd__mux2_1 _06679_ (.A0(_00809_),
    .A1(\Qset[0][4] ),
    .S(_00687_),
    .X(_00810_));
 sky130_fd_sc_hd__clkbuf_1 _06680_ (.A(_00810_),
    .X(_00028_));
 sky130_fd_sc_hd__inv_2 _06681_ (.A(\result_reg_mac[5] ),
    .Y(_00811_));
 sky130_fd_sc_hd__inv_2 _06682_ (.A(\result_reg_add[5] ),
    .Y(_00812_));
 sky130_fd_sc_hd__a21oi_1 _06683_ (.A1(_00541_),
    .A2(_00812_),
    .B1(_00535_),
    .Y(_00813_));
 sky130_fd_sc_hd__o21ai_1 _06684_ (.A1(\result_reg_sub[5] ),
    .A2(_00541_),
    .B1(_00813_),
    .Y(_00814_));
 sky130_fd_sc_hd__inv_2 _06685_ (.A(\result_reg_mul[5] ),
    .Y(_00815_));
 sky130_fd_sc_hd__or2_1 _06686_ (.A(_00815_),
    .B(_00745_),
    .X(_00816_));
 sky130_fd_sc_hd__o21ai_1 _06687_ (.A1(\result_reg_and[5] ),
    .A2(_00562_),
    .B1(_00709_),
    .Y(_00817_));
 sky130_fd_sc_hd__a31o_1 _06688_ (.A1(_00814_),
    .A2(_00562_),
    .A3(_00816_),
    .B1(_00817_),
    .X(_00818_));
 sky130_fd_sc_hd__nand2_1 _06689_ (.A(_00714_),
    .B(\result_reg_or[5] ),
    .Y(_00819_));
 sky130_fd_sc_hd__buf_6 _06690_ (.A(_00710_),
    .X(_00820_));
 sky130_fd_sc_hd__or3_1 _06691_ (.A(CMD_set),
    .B(_00697_),
    .C(_00593_),
    .X(_00821_));
 sky130_fd_sc_hd__or4_1 _06692_ (.A(CMD_not),
    .B(_00545_),
    .C(CMD_and),
    .D(_00821_),
    .X(_00822_));
 sky130_fd_sc_hd__or4_1 _06693_ (.A(\shift.left ),
    .B(CMD_logic_shift_right),
    .C(_00820_),
    .D(_00822_),
    .X(_00823_));
 sky130_fd_sc_hd__or3_1 _06694_ (.A(_00557_),
    .B(_00631_),
    .C(_00823_),
    .X(_00824_));
 sky130_fd_sc_hd__nand2_1 _06695_ (.A(_00592_),
    .B(CMD_set),
    .Y(_00825_));
 sky130_fd_sc_hd__or4_1 _06696_ (.A(CMD_not),
    .B(_00545_),
    .C(CMD_and),
    .D(_00825_),
    .X(_00826_));
 sky130_fd_sc_hd__or4_1 _06697_ (.A(\shift.left ),
    .B(CMD_logic_shift_right),
    .C(_00820_),
    .D(_00826_),
    .X(_00827_));
 sky130_fd_sc_hd__or4_1 _06698_ (.A(_00557_),
    .B(_00631_),
    .C(_00634_),
    .D(_00827_),
    .X(_00828_));
 sky130_fd_sc_hd__inv_2 _06699_ (.A(_00574_),
    .Y(_00829_));
 sky130_fd_sc_hd__or4_1 _06700_ (.A(_00528_),
    .B(_00631_),
    .C(_00634_),
    .D(_00829_),
    .X(_00830_));
 sky130_fd_sc_hd__clkbuf_4 _06701_ (.A(_00536_),
    .X(_00831_));
 sky130_fd_sc_hd__buf_4 _06702_ (.A(_00831_),
    .X(_00832_));
 sky130_fd_sc_hd__inv_2 _06703_ (.A(CMD_addition),
    .Y(_00833_));
 sky130_fd_sc_hd__a2111o_1 _06704_ (.A1(_00832_),
    .A2(_00833_),
    .B1(_06264_),
    .C1(_00635_),
    .D1(_00829_),
    .X(_00834_));
 sky130_fd_sc_hd__o2111ai_4 _06705_ (.A1(_00635_),
    .A2(_00824_),
    .B1(_00828_),
    .C1(_00830_),
    .D1(_00834_),
    .Y(_00835_));
 sky130_fd_sc_hd__a21o_1 _06706_ (.A1(_00818_),
    .A2(_00819_),
    .B1(_00835_),
    .X(_00836_));
 sky130_fd_sc_hd__o211a_1 _06707_ (.A1(_00829_),
    .A2(_00566_),
    .B1(_00732_),
    .C1(_00699_),
    .X(_00837_));
 sky130_fd_sc_hd__and3_1 _06708_ (.A(_00837_),
    .B(_00730_),
    .C(_00607_),
    .X(_00838_));
 sky130_fd_sc_hd__inv_2 _06709_ (.A(_00838_),
    .Y(_00839_));
 sky130_fd_sc_hd__inv_2 _06710_ (.A(\result_reg_set[5] ),
    .Y(_00840_));
 sky130_fd_sc_hd__inv_2 _06711_ (.A(\result_reg_sub[5] ),
    .Y(_00841_));
 sky130_fd_sc_hd__mux2_1 _06712_ (.A0(_00841_),
    .A1(_00812_),
    .S(_00611_),
    .X(_00842_));
 sky130_fd_sc_hd__mux2_1 _06713_ (.A0(_00815_),
    .A1(_00842_),
    .S(_00613_),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_1 _06714_ (.A0(_00840_),
    .A1(_00843_),
    .S(_00608_),
    .X(_00844_));
 sky130_fd_sc_hd__nand2_1 _06715_ (.A(_00844_),
    .B(_00735_),
    .Y(_00845_));
 sky130_fd_sc_hd__o211a_1 _06716_ (.A1(net12),
    .A2(_00735_),
    .B1(_00839_),
    .C1(_00845_),
    .X(_00846_));
 sky130_fd_sc_hd__nor2_1 _06717_ (.A(_00650_),
    .B(_00846_),
    .Y(_00847_));
 sky130_fd_sc_hd__a221o_1 _06718_ (.A1(_00811_),
    .A2(_00695_),
    .B1(_00836_),
    .B2(_00847_),
    .C1(_00644_),
    .X(_00848_));
 sky130_fd_sc_hd__inv_2 _06719_ (.A(\result_reg_not[5] ),
    .Y(_00849_));
 sky130_fd_sc_hd__inv_2 _06720_ (.A(\result_reg_Lshift[5] ),
    .Y(_00850_));
 sky130_fd_sc_hd__nand2_1 _06721_ (.A(_00754_),
    .B(_00850_),
    .Y(_00851_));
 sky130_fd_sc_hd__o21ai_1 _06722_ (.A1(\result_reg_Rshift[5] ),
    .A2(_00753_),
    .B1(_00851_),
    .Y(_00852_));
 sky130_fd_sc_hd__a221o_2 _06723_ (.A1(_00849_),
    .A2(_00655_),
    .B1(_00657_),
    .B2(_00852_),
    .C1(_00666_),
    .X(_00853_));
 sky130_fd_sc_hd__nand2_4 _06724_ (.A(_00848_),
    .B(_00853_),
    .Y(_00854_));
 sky130_fd_sc_hd__mux2_1 _06725_ (.A0(_00854_),
    .A1(\Qset[0][5] ),
    .S(_00687_),
    .X(_00855_));
 sky130_fd_sc_hd__clkbuf_1 _06726_ (.A(_00855_),
    .X(_00029_));
 sky130_fd_sc_hd__inv_2 _06727_ (.A(\result_reg_mac[6] ),
    .Y(_00856_));
 sky130_fd_sc_hd__inv_2 _06728_ (.A(\result_reg_add[6] ),
    .Y(_00857_));
 sky130_fd_sc_hd__a21oi_1 _06729_ (.A1(_00740_),
    .A2(_00857_),
    .B1(_00535_),
    .Y(_00858_));
 sky130_fd_sc_hd__o21ai_1 _06730_ (.A1(\result_reg_sub[6] ),
    .A2(_00541_),
    .B1(_00858_),
    .Y(_00859_));
 sky130_fd_sc_hd__inv_2 _06731_ (.A(\result_reg_mul[6] ),
    .Y(_00860_));
 sky130_fd_sc_hd__or2_1 _06732_ (.A(_00860_),
    .B(_00745_),
    .X(_00861_));
 sky130_fd_sc_hd__o21ai_1 _06733_ (.A1(\result_reg_and[6] ),
    .A2(_00743_),
    .B1(_00553_),
    .Y(_00862_));
 sky130_fd_sc_hd__a31o_1 _06734_ (.A1(_00859_),
    .A2(_00743_),
    .A3(_00861_),
    .B1(_00862_),
    .X(_00863_));
 sky130_fd_sc_hd__or2b_1 _06735_ (.A(_00553_),
    .B_N(\result_reg_or[6] ),
    .X(_00864_));
 sky130_fd_sc_hd__inv_2 _06736_ (.A(\result_reg_sub[6] ),
    .Y(_00865_));
 sky130_fd_sc_hd__mux2_1 _06737_ (.A0(_00865_),
    .A1(_00857_),
    .S(_00730_),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _06738_ (.A0(_00860_),
    .A1(_00866_),
    .S(_00732_),
    .X(_00867_));
 sky130_fd_sc_hd__nand2_1 _06739_ (.A(_00867_),
    .B(_00615_),
    .Y(_00868_));
 sky130_fd_sc_hd__o211ai_1 _06740_ (.A1(\result_reg_set[6] ),
    .A2(_00615_),
    .B1(_00696_),
    .C1(_00868_),
    .Y(_00869_));
 sky130_fd_sc_hd__a21oi_1 _06741_ (.A1(net13),
    .A2(_00600_),
    .B1(_00739_),
    .Y(_00870_));
 sky130_fd_sc_hd__a32o_1 _06742_ (.A1(_00739_),
    .A2(_00863_),
    .A3(_00864_),
    .B1(_00869_),
    .B2(_00870_),
    .X(_00871_));
 sky130_fd_sc_hd__a221o_1 _06743_ (.A1(_00856_),
    .A2(_00695_),
    .B1(_00871_),
    .B2(_00725_),
    .C1(_00644_),
    .X(_00872_));
 sky130_fd_sc_hd__inv_2 _06744_ (.A(\result_reg_not[6] ),
    .Y(_00873_));
 sky130_fd_sc_hd__inv_2 _06745_ (.A(\result_reg_Lshift[6] ),
    .Y(_00874_));
 sky130_fd_sc_hd__nand2_1 _06746_ (.A(_00754_),
    .B(_00874_),
    .Y(_00875_));
 sky130_fd_sc_hd__o21ai_1 _06747_ (.A1(\result_reg_Rshift[6] ),
    .A2(_00753_),
    .B1(_00875_),
    .Y(_00876_));
 sky130_fd_sc_hd__a221o_1 _06748_ (.A1(_00873_),
    .A2(_00655_),
    .B1(_00657_),
    .B2(_00876_),
    .C1(_00666_),
    .X(_00877_));
 sky130_fd_sc_hd__nand2_4 _06749_ (.A(_00872_),
    .B(_00877_),
    .Y(_00878_));
 sky130_fd_sc_hd__mux2_1 _06750_ (.A0(_00878_),
    .A1(\Qset[0][6] ),
    .S(_00687_),
    .X(_00879_));
 sky130_fd_sc_hd__clkbuf_1 _06751_ (.A(_00879_),
    .X(_00030_));
 sky130_fd_sc_hd__inv_2 _06752_ (.A(\result_reg_mac[7] ),
    .Y(_00880_));
 sky130_fd_sc_hd__inv_2 _06753_ (.A(\result_reg_set[7] ),
    .Y(_00881_));
 sky130_fd_sc_hd__inv_2 _06754_ (.A(\result_reg_mul[7] ),
    .Y(_00882_));
 sky130_fd_sc_hd__inv_2 _06755_ (.A(\result_reg_sub[7] ),
    .Y(_00883_));
 sky130_fd_sc_hd__inv_2 _06756_ (.A(\result_reg_add[7] ),
    .Y(_00884_));
 sky130_fd_sc_hd__mux2_1 _06757_ (.A0(_00883_),
    .A1(_00884_),
    .S(_00730_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _06758_ (.A0(_00882_),
    .A1(_00885_),
    .S(_00732_),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_1 _06759_ (.A0(_00881_),
    .A1(_00886_),
    .S(_00608_),
    .X(_00887_));
 sky130_fd_sc_hd__nand2_1 _06760_ (.A(_00887_),
    .B(_00735_),
    .Y(_00888_));
 sky130_fd_sc_hd__o21ai_1 _06761_ (.A1(net14),
    .A2(_00696_),
    .B1(_00888_),
    .Y(_00889_));
 sky130_fd_sc_hd__inv_2 _06762_ (.A(\result_reg_or[7] ),
    .Y(_00890_));
 sky130_fd_sc_hd__a21oi_1 _06763_ (.A1(_00540_),
    .A2(_00884_),
    .B1(_00534_),
    .Y(_00891_));
 sky130_fd_sc_hd__o21ai_1 _06764_ (.A1(\result_reg_sub[7] ),
    .A2(_00740_),
    .B1(_00891_),
    .Y(_00892_));
 sky130_fd_sc_hd__or2_1 _06765_ (.A(_00882_),
    .B(_00745_),
    .X(_00893_));
 sky130_fd_sc_hd__o21ai_1 _06766_ (.A1(\result_reg_and[7] ),
    .A2(_00561_),
    .B1(_00552_),
    .Y(_00894_));
 sky130_fd_sc_hd__a31o_1 _06767_ (.A1(_00892_),
    .A2(_00743_),
    .A3(_00893_),
    .B1(_00894_),
    .X(_00895_));
 sky130_fd_sc_hd__o211a_1 _06768_ (.A1(_00890_),
    .A2(_00709_),
    .B1(_00603_),
    .C1(_00895_),
    .X(_00896_));
 sky130_fd_sc_hd__a211o_1 _06769_ (.A1(_00889_),
    .A2(_00619_),
    .B1(_00629_),
    .C1(_00896_),
    .X(_00897_));
 sky130_fd_sc_hd__o21a_1 _06770_ (.A1(_00880_),
    .A2(_00725_),
    .B1(_00897_),
    .X(_00898_));
 sky130_fd_sc_hd__inv_2 _06771_ (.A(\result_reg_not[7] ),
    .Y(_00899_));
 sky130_fd_sc_hd__inv_2 _06772_ (.A(\result_reg_Rshift[7] ),
    .Y(_00900_));
 sky130_fd_sc_hd__inv_2 _06773_ (.A(\result_reg_Lshift[7] ),
    .Y(_00901_));
 sky130_fd_sc_hd__mux2_1 _06774_ (.A0(_00900_),
    .A1(_00901_),
    .S(_00643_),
    .X(_00902_));
 sky130_fd_sc_hd__a221o_1 _06775_ (.A1(_00899_),
    .A2(_00655_),
    .B1(_00657_),
    .B2(_00902_),
    .C1(_00666_),
    .X(_00903_));
 sky130_fd_sc_hd__o21ai_4 _06776_ (.A1(_00664_),
    .A2(_00898_),
    .B1(_00903_),
    .Y(_00904_));
 sky130_fd_sc_hd__mux2_1 _06777_ (.A0(_00904_),
    .A1(\Qset[0][7] ),
    .S(_00687_),
    .X(_00905_));
 sky130_fd_sc_hd__clkbuf_1 _06778_ (.A(_00905_),
    .X(_00031_));
 sky130_fd_sc_hd__inv_2 _06779_ (.A(\result_reg_add[8] ),
    .Y(_00906_));
 sky130_fd_sc_hd__a21oi_1 _06780_ (.A1(_00541_),
    .A2(_00906_),
    .B1(_00535_),
    .Y(_00907_));
 sky130_fd_sc_hd__or2_1 _06781_ (.A(\result_reg_sub[8] ),
    .B(_00540_),
    .X(_00908_));
 sky130_fd_sc_hd__a221o_1 _06782_ (.A1(\result_reg_mul[8] ),
    .A2(_00535_),
    .B1(_00907_),
    .B2(_00908_),
    .C1(_00563_),
    .X(_00909_));
 sky130_fd_sc_hd__o221a_1 _06783_ (.A1(\result_reg_or[8] ),
    .A2(_00553_),
    .B1(\result_reg_and[8] ),
    .B2(_00562_),
    .C1(_00603_),
    .X(_00910_));
 sky130_fd_sc_hd__inv_2 _06784_ (.A(\result_reg_mul[8] ),
    .Y(_00911_));
 sky130_fd_sc_hd__inv_2 _06785_ (.A(\result_reg_sub[8] ),
    .Y(_00912_));
 sky130_fd_sc_hd__mux2_1 _06786_ (.A0(_00912_),
    .A1(_00906_),
    .S(_00611_),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _06787_ (.A0(_00911_),
    .A1(_00913_),
    .S(_00613_),
    .X(_00914_));
 sky130_fd_sc_hd__nand2_1 _06788_ (.A(_00914_),
    .B(_00615_),
    .Y(_00915_));
 sky130_fd_sc_hd__o211a_1 _06789_ (.A1(\result_reg_set[8] ),
    .A2(_00608_),
    .B1(_00601_),
    .C1(_00915_),
    .X(_00916_));
 sky130_fd_sc_hd__a21o_1 _06790_ (.A1(net15),
    .A2(_00600_),
    .B1(_00916_),
    .X(_00917_));
 sky130_fd_sc_hd__a221o_1 _06791_ (.A1(_00909_),
    .A2(_00910_),
    .B1(_00917_),
    .B2(_00619_),
    .C1(_00629_),
    .X(_00918_));
 sky130_fd_sc_hd__inv_2 _06792_ (.A(\result_reg_mac[8] ),
    .Y(_00919_));
 sky130_fd_sc_hd__nand2_1 _06793_ (.A(_00695_),
    .B(_00919_),
    .Y(_00920_));
 sky130_fd_sc_hd__inv_2 _06794_ (.A(_00654_),
    .Y(_00921_));
 sky130_fd_sc_hd__inv_2 _06795_ (.A(\result_reg_Rshift[8] ),
    .Y(_00922_));
 sky130_fd_sc_hd__inv_2 _06796_ (.A(\result_reg_Lshift[8] ),
    .Y(_00923_));
 sky130_fd_sc_hd__mux2_1 _06797_ (.A0(_00922_),
    .A1(_00923_),
    .S(_00643_),
    .X(_00924_));
 sky130_fd_sc_hd__nand2_1 _06798_ (.A(_00924_),
    .B(_00656_),
    .Y(_00925_));
 sky130_fd_sc_hd__o211a_1 _06799_ (.A1(\result_reg_not[8] ),
    .A2(_00921_),
    .B1(_00925_),
    .C1(_00664_),
    .X(_00926_));
 sky130_fd_sc_hd__a31o_4 _06800_ (.A1(_00918_),
    .A2(_00645_),
    .A3(_00920_),
    .B1(_00926_),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _06801_ (.A0(_00927_),
    .A1(\Qset[0][8] ),
    .S(_00687_),
    .X(_00928_));
 sky130_fd_sc_hd__clkbuf_1 _06802_ (.A(_00928_),
    .X(_00032_));
 sky130_fd_sc_hd__inv_2 _06803_ (.A(\result_reg_mac[9] ),
    .Y(_00929_));
 sky130_fd_sc_hd__inv_2 _06804_ (.A(\result_reg_set[9] ),
    .Y(_00930_));
 sky130_fd_sc_hd__inv_2 _06805_ (.A(\result_reg_mul[9] ),
    .Y(_00931_));
 sky130_fd_sc_hd__inv_2 _06806_ (.A(\result_reg_sub[9] ),
    .Y(_00932_));
 sky130_fd_sc_hd__inv_2 _06807_ (.A(\result_reg_add[9] ),
    .Y(_00933_));
 sky130_fd_sc_hd__mux2_1 _06808_ (.A0(_00932_),
    .A1(_00933_),
    .S(_00730_),
    .X(_00934_));
 sky130_fd_sc_hd__mux2_1 _06809_ (.A0(_00931_),
    .A1(_00934_),
    .S(_00732_),
    .X(_00935_));
 sky130_fd_sc_hd__mux2_1 _06810_ (.A0(_00930_),
    .A1(_00935_),
    .S(_00608_),
    .X(_00936_));
 sky130_fd_sc_hd__nand2_1 _06811_ (.A(_00936_),
    .B(_00735_),
    .Y(_00937_));
 sky130_fd_sc_hd__o21ai_1 _06812_ (.A1(net16),
    .A2(_00696_),
    .B1(_00937_),
    .Y(_00938_));
 sky130_fd_sc_hd__inv_2 _06813_ (.A(\result_reg_or[9] ),
    .Y(_00939_));
 sky130_fd_sc_hd__a21oi_1 _06814_ (.A1(_00540_),
    .A2(_00933_),
    .B1(_00534_),
    .Y(_00940_));
 sky130_fd_sc_hd__o21ai_1 _06815_ (.A1(\result_reg_sub[9] ),
    .A2(_00740_),
    .B1(_00940_),
    .Y(_00941_));
 sky130_fd_sc_hd__or2_1 _06816_ (.A(_00931_),
    .B(_00744_),
    .X(_00942_));
 sky130_fd_sc_hd__o21ai_1 _06817_ (.A1(\result_reg_and[9] ),
    .A2(_00561_),
    .B1(_00552_),
    .Y(_00943_));
 sky130_fd_sc_hd__a31o_1 _06818_ (.A1(_00941_),
    .A2(_00743_),
    .A3(_00942_),
    .B1(_00943_),
    .X(_00944_));
 sky130_fd_sc_hd__o211a_1 _06819_ (.A1(_00939_),
    .A2(_00709_),
    .B1(_00603_),
    .C1(_00944_),
    .X(_00945_));
 sky130_fd_sc_hd__a211o_1 _06820_ (.A1(_00938_),
    .A2(_00619_),
    .B1(_00629_),
    .C1(_00945_),
    .X(_00946_));
 sky130_fd_sc_hd__o21a_1 _06821_ (.A1(_00929_),
    .A2(_00725_),
    .B1(_00946_),
    .X(_00947_));
 sky130_fd_sc_hd__inv_2 _06822_ (.A(\result_reg_not[9] ),
    .Y(_00948_));
 sky130_fd_sc_hd__inv_2 _06823_ (.A(\result_reg_Lshift[9] ),
    .Y(_00949_));
 sky130_fd_sc_hd__nand2_1 _06824_ (.A(_00754_),
    .B(_00949_),
    .Y(_00950_));
 sky130_fd_sc_hd__o21ai_1 _06825_ (.A1(\result_reg_Rshift[9] ),
    .A2(_00753_),
    .B1(_00950_),
    .Y(_00951_));
 sky130_fd_sc_hd__a221o_1 _06826_ (.A1(_00948_),
    .A2(_00655_),
    .B1(_00657_),
    .B2(_00951_),
    .C1(_00666_),
    .X(_00952_));
 sky130_fd_sc_hd__o21ai_4 _06827_ (.A1(_00664_),
    .A2(_00947_),
    .B1(_00952_),
    .Y(_00953_));
 sky130_fd_sc_hd__mux2_1 _06828_ (.A0(_00953_),
    .A1(\Qset[0][9] ),
    .S(_00687_),
    .X(_00954_));
 sky130_fd_sc_hd__clkbuf_1 _06829_ (.A(_00954_),
    .X(_00033_));
 sky130_fd_sc_hd__inv_2 _06830_ (.A(\result_reg_mac[10] ),
    .Y(_00955_));
 sky130_fd_sc_hd__inv_2 _06831_ (.A(\result_reg_set[10] ),
    .Y(_00956_));
 sky130_fd_sc_hd__inv_2 _06832_ (.A(\result_reg_mul[10] ),
    .Y(_00957_));
 sky130_fd_sc_hd__inv_2 _06833_ (.A(\result_reg_sub[10] ),
    .Y(_00958_));
 sky130_fd_sc_hd__inv_2 _06834_ (.A(\result_reg_add[10] ),
    .Y(_00959_));
 sky130_fd_sc_hd__mux2_1 _06835_ (.A0(_00958_),
    .A1(_00959_),
    .S(_00730_),
    .X(_00960_));
 sky130_fd_sc_hd__mux2_1 _06836_ (.A0(_00957_),
    .A1(_00960_),
    .S(_00732_),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_1 _06837_ (.A0(_00956_),
    .A1(_00961_),
    .S(_00608_),
    .X(_00962_));
 sky130_fd_sc_hd__nand2_1 _06838_ (.A(_00962_),
    .B(_00735_),
    .Y(_00963_));
 sky130_fd_sc_hd__o21ai_1 _06839_ (.A1(net2),
    .A2(_00696_),
    .B1(_00963_),
    .Y(_00964_));
 sky130_fd_sc_hd__inv_2 _06840_ (.A(\result_reg_or[10] ),
    .Y(_00965_));
 sky130_fd_sc_hd__a21oi_1 _06841_ (.A1(_00540_),
    .A2(_00959_),
    .B1(_00534_),
    .Y(_00966_));
 sky130_fd_sc_hd__o21ai_1 _06842_ (.A1(\result_reg_sub[10] ),
    .A2(_00740_),
    .B1(_00966_),
    .Y(_00967_));
 sky130_fd_sc_hd__or2_1 _06843_ (.A(_00957_),
    .B(_00744_),
    .X(_00968_));
 sky130_fd_sc_hd__o21ai_1 _06844_ (.A1(\result_reg_and[10] ),
    .A2(_00561_),
    .B1(_00552_),
    .Y(_00969_));
 sky130_fd_sc_hd__a31o_1 _06845_ (.A1(_00967_),
    .A2(_00743_),
    .A3(_00968_),
    .B1(_00969_),
    .X(_00970_));
 sky130_fd_sc_hd__o211a_1 _06846_ (.A1(_00965_),
    .A2(_00709_),
    .B1(_00603_),
    .C1(_00970_),
    .X(_00971_));
 sky130_fd_sc_hd__a211o_1 _06847_ (.A1(_00964_),
    .A2(_00619_),
    .B1(_00629_),
    .C1(_00971_),
    .X(_00972_));
 sky130_fd_sc_hd__o21a_1 _06848_ (.A1(_00955_),
    .A2(_00725_),
    .B1(_00972_),
    .X(_00973_));
 sky130_fd_sc_hd__inv_2 _06849_ (.A(\result_reg_not[10] ),
    .Y(_00974_));
 sky130_fd_sc_hd__inv_2 _06850_ (.A(\result_reg_Lshift[10] ),
    .Y(_00975_));
 sky130_fd_sc_hd__nand2_1 _06851_ (.A(_00754_),
    .B(_00975_),
    .Y(_00976_));
 sky130_fd_sc_hd__o21ai_1 _06852_ (.A1(\result_reg_Rshift[10] ),
    .A2(_00753_),
    .B1(_00976_),
    .Y(_00977_));
 sky130_fd_sc_hd__a221o_1 _06853_ (.A1(_00974_),
    .A2(_00655_),
    .B1(_00657_),
    .B2(_00977_),
    .C1(_00666_),
    .X(_00978_));
 sky130_fd_sc_hd__o21ai_4 _06854_ (.A1(_00664_),
    .A2(_00973_),
    .B1(_00978_),
    .Y(_00979_));
 sky130_fd_sc_hd__mux2_1 _06855_ (.A0(_00979_),
    .A1(\Qset[0][10] ),
    .S(_00686_),
    .X(_00980_));
 sky130_fd_sc_hd__clkbuf_1 _06856_ (.A(_00980_),
    .X(_00034_));
 sky130_fd_sc_hd__inv_2 _06857_ (.A(\result_reg_mac[11] ),
    .Y(_00981_));
 sky130_fd_sc_hd__inv_2 _06858_ (.A(\result_reg_add[11] ),
    .Y(_00982_));
 sky130_fd_sc_hd__a21oi_1 _06859_ (.A1(_00740_),
    .A2(_00982_),
    .B1(_00535_),
    .Y(_00983_));
 sky130_fd_sc_hd__o21ai_1 _06860_ (.A1(\result_reg_sub[11] ),
    .A2(_00541_),
    .B1(_00983_),
    .Y(_00984_));
 sky130_fd_sc_hd__inv_2 _06861_ (.A(\result_reg_mul[11] ),
    .Y(_00985_));
 sky130_fd_sc_hd__or2_1 _06862_ (.A(_00985_),
    .B(_00745_),
    .X(_00986_));
 sky130_fd_sc_hd__o21ai_1 _06863_ (.A1(\result_reg_and[11] ),
    .A2(_00561_),
    .B1(_00553_),
    .Y(_00987_));
 sky130_fd_sc_hd__a31o_1 _06864_ (.A1(_00984_),
    .A2(_00743_),
    .A3(_00986_),
    .B1(_00987_),
    .X(_00988_));
 sky130_fd_sc_hd__inv_2 _06865_ (.A(\result_reg_or[11] ),
    .Y(_00989_));
 sky130_fd_sc_hd__or2_1 _06866_ (.A(_00989_),
    .B(_00553_),
    .X(_00990_));
 sky130_fd_sc_hd__inv_2 _06867_ (.A(\result_reg_sub[11] ),
    .Y(_00991_));
 sky130_fd_sc_hd__mux2_1 _06868_ (.A0(_00991_),
    .A1(_00982_),
    .S(_00730_),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_1 _06869_ (.A0(_00985_),
    .A1(_00992_),
    .S(_00732_),
    .X(_00993_));
 sky130_fd_sc_hd__nand2_1 _06870_ (.A(_00993_),
    .B(_00615_),
    .Y(_00994_));
 sky130_fd_sc_hd__o211ai_1 _06871_ (.A1(\result_reg_set[11] ),
    .A2(_00615_),
    .B1(_00696_),
    .C1(_00994_),
    .Y(_00995_));
 sky130_fd_sc_hd__a21oi_1 _06872_ (.A1(net3),
    .A2(_00600_),
    .B1(_00739_),
    .Y(_00996_));
 sky130_fd_sc_hd__a32o_1 _06873_ (.A1(_00739_),
    .A2(_00988_),
    .A3(_00990_),
    .B1(_00995_),
    .B2(_00996_),
    .X(_00997_));
 sky130_fd_sc_hd__a221o_1 _06874_ (.A1(_00981_),
    .A2(_00695_),
    .B1(_00997_),
    .B2(_00725_),
    .C1(_00644_),
    .X(_00998_));
 sky130_fd_sc_hd__inv_2 _06875_ (.A(\result_reg_not[11] ),
    .Y(_00999_));
 sky130_fd_sc_hd__inv_2 _06876_ (.A(\result_reg_Lshift[11] ),
    .Y(_01000_));
 sky130_fd_sc_hd__nand2_1 _06877_ (.A(_00754_),
    .B(_01000_),
    .Y(_01001_));
 sky130_fd_sc_hd__o21ai_1 _06878_ (.A1(\result_reg_Rshift[11] ),
    .A2(_00753_),
    .B1(_01001_),
    .Y(_01002_));
 sky130_fd_sc_hd__a221o_1 _06879_ (.A1(_00999_),
    .A2(_00655_),
    .B1(_00657_),
    .B2(_01002_),
    .C1(_00666_),
    .X(_01003_));
 sky130_fd_sc_hd__nand2_2 _06880_ (.A(_00998_),
    .B(_01003_),
    .Y(_01004_));
 sky130_fd_sc_hd__mux2_1 _06881_ (.A0(_01004_),
    .A1(\Qset[0][11] ),
    .S(_00686_),
    .X(_01005_));
 sky130_fd_sc_hd__clkbuf_1 _06882_ (.A(_01005_),
    .X(_00035_));
 sky130_fd_sc_hd__inv_2 _06883_ (.A(\result_reg_mac[12] ),
    .Y(_01006_));
 sky130_fd_sc_hd__inv_2 _06884_ (.A(\result_reg_add[12] ),
    .Y(_01007_));
 sky130_fd_sc_hd__a21oi_1 _06885_ (.A1(_00540_),
    .A2(_01007_),
    .B1(_00534_),
    .Y(_01008_));
 sky130_fd_sc_hd__o21ai_1 _06886_ (.A1(\result_reg_sub[12] ),
    .A2(_00541_),
    .B1(_01008_),
    .Y(_01009_));
 sky130_fd_sc_hd__inv_2 _06887_ (.A(\result_reg_mul[12] ),
    .Y(_01010_));
 sky130_fd_sc_hd__or2_1 _06888_ (.A(_01010_),
    .B(_00745_),
    .X(_01011_));
 sky130_fd_sc_hd__o21ai_1 _06889_ (.A1(\result_reg_and[12] ),
    .A2(_00561_),
    .B1(_00552_),
    .Y(_01012_));
 sky130_fd_sc_hd__a31o_1 _06890_ (.A1(_01009_),
    .A2(_00743_),
    .A3(_01011_),
    .B1(_01012_),
    .X(_01013_));
 sky130_fd_sc_hd__inv_2 _06891_ (.A(\result_reg_or[12] ),
    .Y(_01014_));
 sky130_fd_sc_hd__or2_1 _06892_ (.A(_01014_),
    .B(_00553_),
    .X(_01015_));
 sky130_fd_sc_hd__inv_2 _06893_ (.A(\result_reg_sub[12] ),
    .Y(_01016_));
 sky130_fd_sc_hd__mux2_1 _06894_ (.A0(_01016_),
    .A1(_01007_),
    .S(_00730_),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_1 _06895_ (.A0(_01010_),
    .A1(_01017_),
    .S(_00732_),
    .X(_01018_));
 sky130_fd_sc_hd__nand2_1 _06896_ (.A(_01018_),
    .B(_00615_),
    .Y(_01019_));
 sky130_fd_sc_hd__o211ai_1 _06897_ (.A1(\result_reg_set[12] ),
    .A2(_00615_),
    .B1(_00696_),
    .C1(_01019_),
    .Y(_01020_));
 sky130_fd_sc_hd__a21oi_1 _06898_ (.A1(net4),
    .A2(_00600_),
    .B1(_00739_),
    .Y(_01021_));
 sky130_fd_sc_hd__a32o_1 _06899_ (.A1(_00739_),
    .A2(_01013_),
    .A3(_01015_),
    .B1(_01020_),
    .B2(_01021_),
    .X(_01022_));
 sky130_fd_sc_hd__a221o_1 _06900_ (.A1(_01006_),
    .A2(_00695_),
    .B1(_01022_),
    .B2(_00725_),
    .C1(_00644_),
    .X(_01023_));
 sky130_fd_sc_hd__inv_2 _06901_ (.A(\result_reg_not[12] ),
    .Y(_01024_));
 sky130_fd_sc_hd__inv_2 _06902_ (.A(\result_reg_Lshift[12] ),
    .Y(_01025_));
 sky130_fd_sc_hd__nand2_1 _06903_ (.A(_00754_),
    .B(_01025_),
    .Y(_01026_));
 sky130_fd_sc_hd__o21ai_1 _06904_ (.A1(\result_reg_Rshift[12] ),
    .A2(_00753_),
    .B1(_01026_),
    .Y(_01027_));
 sky130_fd_sc_hd__a221o_1 _06905_ (.A1(_01024_),
    .A2(_00654_),
    .B1(_00656_),
    .B2(_01027_),
    .C1(_00665_),
    .X(_01028_));
 sky130_fd_sc_hd__nand2_2 _06906_ (.A(_01023_),
    .B(_01028_),
    .Y(_01029_));
 sky130_fd_sc_hd__mux2_1 _06907_ (.A0(_01029_),
    .A1(\Qset[0][12] ),
    .S(_00686_),
    .X(_01030_));
 sky130_fd_sc_hd__clkbuf_1 _06908_ (.A(_01030_),
    .X(_00036_));
 sky130_fd_sc_hd__inv_2 _06909_ (.A(\result_reg_mac[13] ),
    .Y(_01031_));
 sky130_fd_sc_hd__inv_2 _06910_ (.A(net5),
    .Y(_01032_));
 sky130_fd_sc_hd__inv_2 _06911_ (.A(\result_reg_set[13] ),
    .Y(_01033_));
 sky130_fd_sc_hd__inv_2 _06912_ (.A(\result_reg_mul[13] ),
    .Y(_01034_));
 sky130_fd_sc_hd__inv_2 _06913_ (.A(\result_reg_sub[13] ),
    .Y(_01035_));
 sky130_fd_sc_hd__inv_2 _06914_ (.A(\result_reg_add[13] ),
    .Y(_01036_));
 sky130_fd_sc_hd__mux2_1 _06915_ (.A0(_01035_),
    .A1(_01036_),
    .S(_00611_),
    .X(_01037_));
 sky130_fd_sc_hd__mux2_1 _06916_ (.A0(_01034_),
    .A1(_01037_),
    .S(_00613_),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_1 _06917_ (.A0(_01033_),
    .A1(_01038_),
    .S(_00607_),
    .X(_01039_));
 sky130_fd_sc_hd__a22o_1 _06918_ (.A1(_01032_),
    .A2(_00600_),
    .B1(_01039_),
    .B2(_00699_),
    .X(_01040_));
 sky130_fd_sc_hd__inv_2 _06919_ (.A(\result_reg_or[13] ),
    .Y(_01041_));
 sky130_fd_sc_hd__inv_2 _06920_ (.A(\result_reg_and[13] ),
    .Y(_01042_));
 sky130_fd_sc_hd__mux2_1 _06921_ (.A0(_01035_),
    .A1(_01036_),
    .S(_00539_),
    .X(_01043_));
 sky130_fd_sc_hd__mux2_1 _06922_ (.A0(_01043_),
    .A1(_01034_),
    .S(_00534_),
    .X(_01044_));
 sky130_fd_sc_hd__mux2_1 _06923_ (.A0(_01042_),
    .A1(_01044_),
    .S(_00561_),
    .X(_01045_));
 sky130_fd_sc_hd__o221a_1 _06924_ (.A1(_01041_),
    .A2(_00709_),
    .B1(_00714_),
    .B2(_01045_),
    .C1(_00603_),
    .X(_01046_));
 sky130_fd_sc_hd__a21o_1 _06925_ (.A1(_01040_),
    .A2(_00619_),
    .B1(_01046_),
    .X(_01047_));
 sky130_fd_sc_hd__a221o_1 _06926_ (.A1(_01031_),
    .A2(_00695_),
    .B1(_01047_),
    .B2(_00725_),
    .C1(_00644_),
    .X(_01048_));
 sky130_fd_sc_hd__inv_2 _06927_ (.A(\result_reg_not[13] ),
    .Y(_01049_));
 sky130_fd_sc_hd__inv_2 _06928_ (.A(\result_reg_Lshift[13] ),
    .Y(_01050_));
 sky130_fd_sc_hd__nand2_1 _06929_ (.A(_00754_),
    .B(_01050_),
    .Y(_01051_));
 sky130_fd_sc_hd__o21ai_1 _06930_ (.A1(\result_reg_Rshift[13] ),
    .A2(_00753_),
    .B1(_01051_),
    .Y(_01052_));
 sky130_fd_sc_hd__a221o_1 _06931_ (.A1(_01049_),
    .A2(_00654_),
    .B1(_00656_),
    .B2(_01052_),
    .C1(_00665_),
    .X(_01053_));
 sky130_fd_sc_hd__nand2_2 _06932_ (.A(_01048_),
    .B(_01053_),
    .Y(_01054_));
 sky130_fd_sc_hd__mux2_1 _06933_ (.A0(_01054_),
    .A1(\Qset[0][13] ),
    .S(_00686_),
    .X(_01055_));
 sky130_fd_sc_hd__clkbuf_1 _06934_ (.A(_01055_),
    .X(_00037_));
 sky130_fd_sc_hd__inv_2 _06935_ (.A(\result_reg_mac[14] ),
    .Y(_01056_));
 sky130_fd_sc_hd__inv_2 _06936_ (.A(\result_reg_add[14] ),
    .Y(_01057_));
 sky130_fd_sc_hd__a21oi_1 _06937_ (.A1(_00740_),
    .A2(_01057_),
    .B1(_00535_),
    .Y(_01058_));
 sky130_fd_sc_hd__o21ai_2 _06938_ (.A1(\result_reg_sub[14] ),
    .A2(_00541_),
    .B1(_01058_),
    .Y(_01059_));
 sky130_fd_sc_hd__inv_2 _06939_ (.A(\result_reg_mul[14] ),
    .Y(_01060_));
 sky130_fd_sc_hd__or2_1 _06940_ (.A(_01060_),
    .B(_00745_),
    .X(_01061_));
 sky130_fd_sc_hd__o21ai_1 _06941_ (.A1(\result_reg_and[14] ),
    .A2(_00562_),
    .B1(_00709_),
    .Y(_01062_));
 sky130_fd_sc_hd__a31o_1 _06942_ (.A1(_01059_),
    .A2(_00562_),
    .A3(_01061_),
    .B1(_01062_),
    .X(_01063_));
 sky130_fd_sc_hd__nand2_1 _06943_ (.A(_00714_),
    .B(\result_reg_or[14] ),
    .Y(_01064_));
 sky130_fd_sc_hd__a21o_1 _06944_ (.A1(_01063_),
    .A2(_01064_),
    .B1(_00835_),
    .X(_01065_));
 sky130_fd_sc_hd__inv_2 _06945_ (.A(\result_reg_set[14] ),
    .Y(_01066_));
 sky130_fd_sc_hd__inv_2 _06946_ (.A(\result_reg_sub[14] ),
    .Y(_01067_));
 sky130_fd_sc_hd__mux2_1 _06947_ (.A0(_01067_),
    .A1(_01057_),
    .S(_00611_),
    .X(_01068_));
 sky130_fd_sc_hd__mux2_1 _06948_ (.A0(_01060_),
    .A1(_01068_),
    .S(_00613_),
    .X(_01069_));
 sky130_fd_sc_hd__mux2_1 _06949_ (.A0(_01066_),
    .A1(_01069_),
    .S(_00608_),
    .X(_01070_));
 sky130_fd_sc_hd__nand2_1 _06950_ (.A(_01070_),
    .B(_00735_),
    .Y(_01071_));
 sky130_fd_sc_hd__o211a_1 _06951_ (.A1(net6),
    .A2(_00735_),
    .B1(_00839_),
    .C1(_01071_),
    .X(_01072_));
 sky130_fd_sc_hd__nor2_1 _06952_ (.A(_00650_),
    .B(_01072_),
    .Y(_01073_));
 sky130_fd_sc_hd__a221o_1 _06953_ (.A1(_01056_),
    .A2(_00695_),
    .B1(_01065_),
    .B2(_01073_),
    .C1(_00644_),
    .X(_01074_));
 sky130_fd_sc_hd__inv_2 _06954_ (.A(\result_reg_not[14] ),
    .Y(_01075_));
 sky130_fd_sc_hd__inv_2 _06955_ (.A(\result_reg_Lshift[14] ),
    .Y(_01076_));
 sky130_fd_sc_hd__nand2_1 _06956_ (.A(_00754_),
    .B(_01076_),
    .Y(_01077_));
 sky130_fd_sc_hd__o21ai_1 _06957_ (.A1(\result_reg_Rshift[14] ),
    .A2(_00753_),
    .B1(_01077_),
    .Y(_01078_));
 sky130_fd_sc_hd__a221o_1 _06958_ (.A1(_01075_),
    .A2(_00654_),
    .B1(_00656_),
    .B2(_01078_),
    .C1(_00665_),
    .X(_01079_));
 sky130_fd_sc_hd__nand2_1 _06959_ (.A(_01074_),
    .B(_01079_),
    .Y(_01080_));
 sky130_fd_sc_hd__mux2_1 _06960_ (.A0(_01080_),
    .A1(\Qset[0][14] ),
    .S(_00686_),
    .X(_01081_));
 sky130_fd_sc_hd__clkbuf_1 _06961_ (.A(_01081_),
    .X(_00038_));
 sky130_fd_sc_hd__inv_2 _06962_ (.A(\result_reg_mac[15] ),
    .Y(_01082_));
 sky130_fd_sc_hd__inv_2 _06963_ (.A(\result_reg_add[15] ),
    .Y(_01083_));
 sky130_fd_sc_hd__a21oi_1 _06964_ (.A1(_00740_),
    .A2(_01083_),
    .B1(_00535_),
    .Y(_01084_));
 sky130_fd_sc_hd__o21ai_2 _06965_ (.A1(\result_reg_sub[15] ),
    .A2(_00541_),
    .B1(_01084_),
    .Y(_01085_));
 sky130_fd_sc_hd__inv_2 _06966_ (.A(\result_reg_mul[15] ),
    .Y(_01086_));
 sky130_fd_sc_hd__or2_1 _06967_ (.A(_01086_),
    .B(_00745_),
    .X(_01087_));
 sky130_fd_sc_hd__o21ai_1 _06968_ (.A1(\result_reg_and[15] ),
    .A2(_00562_),
    .B1(_00709_),
    .Y(_01088_));
 sky130_fd_sc_hd__a31o_1 _06969_ (.A1(_01085_),
    .A2(_00562_),
    .A3(_01087_),
    .B1(_01088_),
    .X(_01089_));
 sky130_fd_sc_hd__nand2_1 _06970_ (.A(_00714_),
    .B(\result_reg_or[15] ),
    .Y(_01090_));
 sky130_fd_sc_hd__a21o_1 _06971_ (.A1(_01089_),
    .A2(_01090_),
    .B1(_00835_),
    .X(_01091_));
 sky130_fd_sc_hd__inv_2 _06972_ (.A(\result_reg_set[15] ),
    .Y(_01092_));
 sky130_fd_sc_hd__inv_2 _06973_ (.A(\result_reg_sub[15] ),
    .Y(_01093_));
 sky130_fd_sc_hd__mux2_1 _06974_ (.A0(_01093_),
    .A1(_01083_),
    .S(_00611_),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_1 _06975_ (.A0(_01086_),
    .A1(_01094_),
    .S(_00613_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _06976_ (.A0(_01092_),
    .A1(_01095_),
    .S(_00608_),
    .X(_01096_));
 sky130_fd_sc_hd__nand2_1 _06977_ (.A(_01096_),
    .B(_00735_),
    .Y(_01097_));
 sky130_fd_sc_hd__o211a_1 _06978_ (.A1(net7),
    .A2(_00699_),
    .B1(_00839_),
    .C1(_01097_),
    .X(_01098_));
 sky130_fd_sc_hd__nor2_1 _06979_ (.A(_00650_),
    .B(_01098_),
    .Y(_01099_));
 sky130_fd_sc_hd__a221o_1 _06980_ (.A1(_01082_),
    .A2(_00695_),
    .B1(_01091_),
    .B2(_01099_),
    .C1(_00644_),
    .X(_01100_));
 sky130_fd_sc_hd__inv_2 _06981_ (.A(\result_reg_not[15] ),
    .Y(_01101_));
 sky130_fd_sc_hd__inv_2 _06982_ (.A(\result_reg_Rshift[15] ),
    .Y(_01102_));
 sky130_fd_sc_hd__inv_2 _06983_ (.A(\result_reg_Lshift[15] ),
    .Y(_01103_));
 sky130_fd_sc_hd__mux2_1 _06984_ (.A0(_01102_),
    .A1(_01103_),
    .S(_00643_),
    .X(_01104_));
 sky130_fd_sc_hd__a221o_1 _06985_ (.A1(_01101_),
    .A2(_00654_),
    .B1(_00656_),
    .B2(_01104_),
    .C1(_00665_),
    .X(_01105_));
 sky130_fd_sc_hd__nand2_1 _06986_ (.A(_01100_),
    .B(_01105_),
    .Y(_01106_));
 sky130_fd_sc_hd__mux2_1 _06987_ (.A0(_01106_),
    .A1(\Qset[0][15] ),
    .S(_00686_),
    .X(_01107_));
 sky130_fd_sc_hd__clkbuf_1 _06988_ (.A(_01107_),
    .X(_00039_));
 sky130_fd_sc_hd__nand2_4 _06989_ (.A(_00679_),
    .B(_00684_),
    .Y(_01108_));
 sky130_fd_sc_hd__clkbuf_8 _06990_ (.A(_01108_),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _06991_ (.A0(_00668_),
    .A1(\Qset[1][0] ),
    .S(_01109_),
    .X(_01110_));
 sky130_fd_sc_hd__clkbuf_1 _06992_ (.A(_01110_),
    .X(_00040_));
 sky130_fd_sc_hd__mux2_1 _06993_ (.A0(_00722_),
    .A1(\Qset[1][1] ),
    .S(_01109_),
    .X(_01111_));
 sky130_fd_sc_hd__clkbuf_1 _06994_ (.A(_01111_),
    .X(_00041_));
 sky130_fd_sc_hd__mux2_1 _06995_ (.A0(_00759_),
    .A1(\Qset[1][2] ),
    .S(_01109_),
    .X(_01112_));
 sky130_fd_sc_hd__clkbuf_1 _06996_ (.A(_01112_),
    .X(_00042_));
 sky130_fd_sc_hd__mux2_1 _06997_ (.A0(_00783_),
    .A1(\Qset[1][3] ),
    .S(_01109_),
    .X(_01113_));
 sky130_fd_sc_hd__clkbuf_1 _06998_ (.A(_01113_),
    .X(_00043_));
 sky130_fd_sc_hd__mux2_1 _06999_ (.A0(_00809_),
    .A1(\Qset[1][4] ),
    .S(_01109_),
    .X(_01114_));
 sky130_fd_sc_hd__clkbuf_1 _07000_ (.A(_01114_),
    .X(_00044_));
 sky130_fd_sc_hd__mux2_1 _07001_ (.A0(_00854_),
    .A1(\Qset[1][5] ),
    .S(_01109_),
    .X(_01115_));
 sky130_fd_sc_hd__clkbuf_1 _07002_ (.A(_01115_),
    .X(_00045_));
 sky130_fd_sc_hd__mux2_1 _07003_ (.A0(_00878_),
    .A1(\Qset[1][6] ),
    .S(_01109_),
    .X(_01116_));
 sky130_fd_sc_hd__clkbuf_1 _07004_ (.A(_01116_),
    .X(_00046_));
 sky130_fd_sc_hd__mux2_1 _07005_ (.A0(_00904_),
    .A1(\Qset[1][7] ),
    .S(_01109_),
    .X(_01117_));
 sky130_fd_sc_hd__clkbuf_1 _07006_ (.A(_01117_),
    .X(_00047_));
 sky130_fd_sc_hd__mux2_1 _07007_ (.A0(_00927_),
    .A1(\Qset[1][8] ),
    .S(_01109_),
    .X(_01118_));
 sky130_fd_sc_hd__clkbuf_1 _07008_ (.A(_01118_),
    .X(_00048_));
 sky130_fd_sc_hd__mux2_1 _07009_ (.A0(_00953_),
    .A1(\Qset[1][9] ),
    .S(_01109_),
    .X(_01119_));
 sky130_fd_sc_hd__clkbuf_1 _07010_ (.A(_01119_),
    .X(_00049_));
 sky130_fd_sc_hd__mux2_1 _07011_ (.A0(_00979_),
    .A1(\Qset[1][10] ),
    .S(_01108_),
    .X(_01120_));
 sky130_fd_sc_hd__clkbuf_1 _07012_ (.A(_01120_),
    .X(_00050_));
 sky130_fd_sc_hd__mux2_1 _07013_ (.A0(_01004_),
    .A1(\Qset[1][11] ),
    .S(_01108_),
    .X(_01121_));
 sky130_fd_sc_hd__clkbuf_1 _07014_ (.A(_01121_),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _07015_ (.A0(_01029_),
    .A1(\Qset[1][12] ),
    .S(_01108_),
    .X(_01122_));
 sky130_fd_sc_hd__clkbuf_1 _07016_ (.A(_01122_),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _07017_ (.A0(_01054_),
    .A1(\Qset[1][13] ),
    .S(_01108_),
    .X(_01123_));
 sky130_fd_sc_hd__clkbuf_1 _07018_ (.A(_01123_),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _07019_ (.A0(_01080_),
    .A1(\Qset[1][14] ),
    .S(_01108_),
    .X(_01124_));
 sky130_fd_sc_hd__clkbuf_1 _07020_ (.A(_01124_),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _07021_ (.A0(_01106_),
    .A1(\Qset[1][15] ),
    .S(_01108_),
    .X(_01125_));
 sky130_fd_sc_hd__clkbuf_1 _07022_ (.A(_01125_),
    .X(_00055_));
 sky130_fd_sc_hd__or2b_1 _07023_ (.A(_00675_),
    .B_N(_00677_),
    .X(_01126_));
 sky130_fd_sc_hd__or2_1 _07024_ (.A(_00684_),
    .B(_01126_),
    .X(_01127_));
 sky130_fd_sc_hd__clkbuf_4 _07025_ (.A(_01127_),
    .X(_01128_));
 sky130_fd_sc_hd__clkbuf_8 _07026_ (.A(_01128_),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_1 _07027_ (.A0(_00668_),
    .A1(\Qset[2][0] ),
    .S(_01129_),
    .X(_01130_));
 sky130_fd_sc_hd__clkbuf_1 _07028_ (.A(_01130_),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _07029_ (.A0(_00722_),
    .A1(\Qset[2][1] ),
    .S(_01129_),
    .X(_01131_));
 sky130_fd_sc_hd__clkbuf_1 _07030_ (.A(_01131_),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _07031_ (.A0(_00759_),
    .A1(\Qset[2][2] ),
    .S(_01129_),
    .X(_01132_));
 sky130_fd_sc_hd__clkbuf_1 _07032_ (.A(_01132_),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _07033_ (.A0(_00783_),
    .A1(\Qset[2][3] ),
    .S(_01129_),
    .X(_01133_));
 sky130_fd_sc_hd__clkbuf_1 _07034_ (.A(_01133_),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _07035_ (.A0(_00809_),
    .A1(\Qset[2][4] ),
    .S(_01129_),
    .X(_01134_));
 sky130_fd_sc_hd__clkbuf_1 _07036_ (.A(_01134_),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _07037_ (.A0(_00854_),
    .A1(\Qset[2][5] ),
    .S(_01129_),
    .X(_01135_));
 sky130_fd_sc_hd__clkbuf_1 _07038_ (.A(_01135_),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _07039_ (.A0(_00878_),
    .A1(\Qset[2][6] ),
    .S(_01129_),
    .X(_01136_));
 sky130_fd_sc_hd__clkbuf_1 _07040_ (.A(_01136_),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _07041_ (.A0(_00904_),
    .A1(\Qset[2][7] ),
    .S(_01129_),
    .X(_01137_));
 sky130_fd_sc_hd__clkbuf_1 _07042_ (.A(_01137_),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_1 _07043_ (.A0(_00927_),
    .A1(\Qset[2][8] ),
    .S(_01129_),
    .X(_01138_));
 sky130_fd_sc_hd__clkbuf_1 _07044_ (.A(_01138_),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _07045_ (.A0(_00953_),
    .A1(\Qset[2][9] ),
    .S(_01129_),
    .X(_01139_));
 sky130_fd_sc_hd__clkbuf_1 _07046_ (.A(_01139_),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _07047_ (.A0(_00979_),
    .A1(\Qset[2][10] ),
    .S(_01128_),
    .X(_01140_));
 sky130_fd_sc_hd__clkbuf_1 _07048_ (.A(_01140_),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _07049_ (.A0(_01004_),
    .A1(\Qset[2][11] ),
    .S(_01128_),
    .X(_01141_));
 sky130_fd_sc_hd__clkbuf_1 _07050_ (.A(_01141_),
    .X(_00067_));
 sky130_fd_sc_hd__mux2_1 _07051_ (.A0(_01029_),
    .A1(\Qset[2][12] ),
    .S(_01128_),
    .X(_01142_));
 sky130_fd_sc_hd__clkbuf_1 _07052_ (.A(_01142_),
    .X(_00068_));
 sky130_fd_sc_hd__mux2_1 _07053_ (.A0(_01054_),
    .A1(\Qset[2][13] ),
    .S(_01128_),
    .X(_01143_));
 sky130_fd_sc_hd__clkbuf_1 _07054_ (.A(_01143_),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _07055_ (.A0(_01080_),
    .A1(\Qset[2][14] ),
    .S(_01128_),
    .X(_01144_));
 sky130_fd_sc_hd__clkbuf_1 _07056_ (.A(_01144_),
    .X(_00070_));
 sky130_fd_sc_hd__mux2_1 _07057_ (.A0(_01106_),
    .A1(\Qset[2][15] ),
    .S(_01128_),
    .X(_01145_));
 sky130_fd_sc_hd__clkbuf_1 _07058_ (.A(_01145_),
    .X(_00071_));
 sky130_fd_sc_hd__clkbuf_4 _07059_ (.A(\current_state[2] ),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _07060_ (.A0(\R0[0] ),
    .A1(net18),
    .S(_01146_),
    .X(_01147_));
 sky130_fd_sc_hd__clkbuf_4 _07061_ (.A(_00472_),
    .X(_01148_));
 sky130_fd_sc_hd__buf_6 _07062_ (.A(_01148_),
    .X(_01149_));
 sky130_fd_sc_hd__and2_1 _07063_ (.A(_01147_),
    .B(_01149_),
    .X(_01150_));
 sky130_fd_sc_hd__clkbuf_1 _07064_ (.A(_01150_),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _07065_ (.A0(\R0[1] ),
    .A1(net19),
    .S(\current_state[2] ),
    .X(_01151_));
 sky130_fd_sc_hd__and2_1 _07066_ (.A(_01151_),
    .B(_01149_),
    .X(_01152_));
 sky130_fd_sc_hd__buf_1 _07067_ (.A(_01152_),
    .X(_00073_));
 sky130_fd_sc_hd__inv_2 _07068_ (.A(_00583_),
    .Y(_01153_));
 sky130_fd_sc_hd__buf_4 _07069_ (.A(_01153_),
    .X(_01154_));
 sky130_fd_sc_hd__buf_4 _07070_ (.A(_01154_),
    .X(_01155_));
 sky130_fd_sc_hd__clkbuf_4 _07071_ (.A(_01155_),
    .X(_01156_));
 sky130_fd_sc_hd__nor2_2 _07072_ (.A(_00589_),
    .B(_01156_),
    .Y(_01157_));
 sky130_fd_sc_hd__buf_4 _07073_ (.A(_01157_),
    .X(_01158_));
 sky130_fd_sc_hd__o311a_4 _07074_ (.A1(_00641_),
    .A2(_00640_),
    .A3(_00654_),
    .B1(_00530_),
    .C1(_01158_),
    .X(_01159_));
 sky130_fd_sc_hd__buf_2 _07075_ (.A(_01159_),
    .X(_01160_));
 sky130_fd_sc_hd__buf_4 _07076_ (.A(_01160_),
    .X(_01161_));
 sky130_fd_sc_hd__inv_2 _07077_ (.A(_01157_),
    .Y(_01162_));
 sky130_fd_sc_hd__nor2_2 _07078_ (.A(_01162_),
    .B(_00531_),
    .Y(_01163_));
 sky130_fd_sc_hd__nand2_4 _07079_ (.A(_01163_),
    .B(_00641_),
    .Y(_01164_));
 sky130_fd_sc_hd__buf_4 _07080_ (.A(_01164_),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _07081_ (.A0(\result_reg_Lshift[0] ),
    .A1(\result_reg_Rshift[0] ),
    .S(_01165_),
    .X(_01166_));
 sky130_fd_sc_hd__nand2_4 _07082_ (.A(_01163_),
    .B(_00654_),
    .Y(_01167_));
 sky130_fd_sc_hd__buf_4 _07083_ (.A(_01167_),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _07084_ (.A0(\result_reg_not[0] ),
    .A1(_01166_),
    .S(_01168_),
    .X(_01169_));
 sky130_fd_sc_hd__inv_2 _07085_ (.A(\result_reg_set[0] ),
    .Y(_01170_));
 sky130_fd_sc_hd__or3_2 _07086_ (.A(_00570_),
    .B(Him),
    .C(_00573_),
    .X(_01171_));
 sky130_fd_sc_hd__inv_2 _07087_ (.A(_01171_),
    .Y(_01172_));
 sky130_fd_sc_hd__nand2_4 _07088_ (.A(_00538_),
    .B(_01172_),
    .Y(_01173_));
 sky130_fd_sc_hd__buf_4 _07089_ (.A(_01173_),
    .X(_01174_));
 sky130_fd_sc_hd__mux2_1 _07090_ (.A0(_00610_),
    .A1(_00542_),
    .S(_01174_),
    .X(_01175_));
 sky130_fd_sc_hd__nand2_4 _07091_ (.A(_01172_),
    .B(_00532_),
    .Y(_01176_));
 sky130_fd_sc_hd__buf_4 _07092_ (.A(_01176_),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _07093_ (.A0(_00609_),
    .A1(_01175_),
    .S(_01177_),
    .X(_01178_));
 sky130_fd_sc_hd__and3_1 _07094_ (.A(_00471_),
    .B(_00558_),
    .C(_01157_),
    .X(_01179_));
 sky130_fd_sc_hd__nor2_1 _07095_ (.A(_00579_),
    .B(_00653_),
    .Y(_01180_));
 sky130_fd_sc_hd__nand2_4 _07096_ (.A(_01179_),
    .B(_01180_),
    .Y(_01181_));
 sky130_fd_sc_hd__clkbuf_4 _07097_ (.A(_01181_),
    .X(_01182_));
 sky130_fd_sc_hd__mux2_1 _07098_ (.A0(_01170_),
    .A1(_01178_),
    .S(_01182_),
    .X(_01183_));
 sky130_fd_sc_hd__nor2_1 _07099_ (.A(_00698_),
    .B(_00653_),
    .Y(_01184_));
 sky130_fd_sc_hd__and3_2 _07100_ (.A(_01179_),
    .B(CMD_load),
    .C(_01184_),
    .X(_01185_));
 sky130_fd_sc_hd__inv_2 _07101_ (.A(_01185_),
    .Y(_01186_));
 sky130_fd_sc_hd__buf_2 _07102_ (.A(_01186_),
    .X(_01187_));
 sky130_fd_sc_hd__nor2_1 _07103_ (.A(_01171_),
    .B(_00568_),
    .Y(_01188_));
 sky130_fd_sc_hd__or3b_1 _07104_ (.A(_01185_),
    .B(_01188_),
    .C_N(_01181_),
    .X(_01189_));
 sky130_fd_sc_hd__clkbuf_4 _07105_ (.A(_01189_),
    .X(_01190_));
 sky130_fd_sc_hd__inv_2 _07106_ (.A(_01190_),
    .Y(_01191_));
 sky130_fd_sc_hd__clkbuf_4 _07107_ (.A(_01191_),
    .X(_01192_));
 sky130_fd_sc_hd__buf_2 _07108_ (.A(_01186_),
    .X(_01193_));
 sky130_fd_sc_hd__nor2_1 _07109_ (.A(net1),
    .B(_01193_),
    .Y(_01194_));
 sky130_fd_sc_hd__a211o_1 _07110_ (.A1(_01183_),
    .A2(_01187_),
    .B1(_01192_),
    .C1(_01194_),
    .X(_01195_));
 sky130_fd_sc_hd__and4_2 _07111_ (.A(_00550_),
    .B(_00471_),
    .C(_00545_),
    .D(_00558_),
    .X(_01196_));
 sky130_fd_sc_hd__inv_2 _07112_ (.A(Oreg2),
    .Y(_01197_));
 sky130_fd_sc_hd__nor2_4 _07113_ (.A(Hreg2),
    .B(_01197_),
    .Y(_01198_));
 sky130_fd_sc_hd__nand2_4 _07114_ (.A(_01196_),
    .B(_01198_),
    .Y(_01199_));
 sky130_fd_sc_hd__clkinv_4 _07115_ (.A(_01198_),
    .Y(_01200_));
 sky130_fd_sc_hd__nor2_1 _07116_ (.A(_01200_),
    .B(_00537_),
    .Y(_01201_));
 sky130_fd_sc_hd__buf_4 _07117_ (.A(_01201_),
    .X(_01202_));
 sky130_fd_sc_hd__mux2_1 _07118_ (.A0(\result_reg_add[0] ),
    .A1(\result_reg_sub[0] ),
    .S(_01202_),
    .X(_01203_));
 sky130_fd_sc_hd__nor2_4 _07119_ (.A(_01200_),
    .B(_00533_),
    .Y(_01204_));
 sky130_fd_sc_hd__mux2_1 _07120_ (.A0(_01203_),
    .A1(\result_reg_mul[0] ),
    .S(_01204_),
    .X(_01205_));
 sky130_fd_sc_hd__nand2_2 _07121_ (.A(_00559_),
    .B(_01198_),
    .Y(_01206_));
 sky130_fd_sc_hd__clkbuf_4 _07122_ (.A(_01206_),
    .X(_01207_));
 sky130_fd_sc_hd__inv_2 _07123_ (.A(_01199_),
    .Y(_01208_));
 sky130_fd_sc_hd__inv_2 _07124_ (.A(\result_reg_and[0] ),
    .Y(_01209_));
 sky130_fd_sc_hd__nor2_1 _07125_ (.A(_01209_),
    .B(_01207_),
    .Y(_01210_));
 sky130_fd_sc_hd__a211o_1 _07126_ (.A1(_01205_),
    .A2(_01207_),
    .B1(_01208_),
    .C1(_01210_),
    .X(_01211_));
 sky130_fd_sc_hd__o211ai_1 _07127_ (.A1(\result_reg_or[0] ),
    .A2(_01199_),
    .B1(_01192_),
    .C1(_01211_),
    .Y(_01212_));
 sky130_fd_sc_hd__or3_1 _07128_ (.A(_00647_),
    .B(_00625_),
    .C(_00627_),
    .X(_01213_));
 sky130_fd_sc_hd__clkbuf_4 _07129_ (.A(_01213_),
    .X(_01214_));
 sky130_fd_sc_hd__clkbuf_4 _07130_ (.A(_01214_),
    .X(_01215_));
 sky130_fd_sc_hd__nor2_1 _07131_ (.A(\result_reg_mac[0] ),
    .B(_01215_),
    .Y(_01216_));
 sky130_fd_sc_hd__a311o_1 _07132_ (.A1(_01195_),
    .A2(_01212_),
    .A3(_01214_),
    .B1(_01160_),
    .C1(_01216_),
    .X(_01217_));
 sky130_fd_sc_hd__a21bo_4 _07133_ (.A1(_01161_),
    .A2(_01169_),
    .B1_N(_01217_),
    .X(_01218_));
 sky130_fd_sc_hd__o21ai_2 _07134_ (.A1(_00661_),
    .A2(_00654_),
    .B1(_01163_),
    .Y(_01219_));
 sky130_fd_sc_hd__inv_2 _07135_ (.A(_01214_),
    .Y(_01220_));
 sky130_fd_sc_hd__nand2_1 _07136_ (.A(_01190_),
    .B(\R0[0] ),
    .Y(_01221_));
 sky130_fd_sc_hd__o21a_1 _07137_ (.A1(_00681_),
    .A2(_01190_),
    .B1(_01221_),
    .X(_01222_));
 sky130_fd_sc_hd__nor2_1 _07138_ (.A(_01220_),
    .B(_01222_),
    .Y(_01223_));
 sky130_fd_sc_hd__a211o_1 _07139_ (.A1(_00498_),
    .A2(_01220_),
    .B1(_01159_),
    .C1(_01223_),
    .X(_01224_));
 sky130_fd_sc_hd__o21ai_4 _07140_ (.A1(\R3[0] ),
    .A2(_01219_),
    .B1(_01224_),
    .Y(_01225_));
 sky130_fd_sc_hd__inv_2 _07141_ (.A(\R1[1] ),
    .Y(_01226_));
 sky130_fd_sc_hd__nor2_1 _07142_ (.A(_01226_),
    .B(_01214_),
    .Y(_01227_));
 sky130_fd_sc_hd__or3_1 _07143_ (.A(CMD_set),
    .B(_00697_),
    .C(_01162_),
    .X(_01228_));
 sky130_fd_sc_hd__or4_1 _07144_ (.A(CMD_not),
    .B(_00545_),
    .C(CMD_and),
    .D(_01228_),
    .X(_01229_));
 sky130_fd_sc_hd__or4_1 _07145_ (.A(\shift.left ),
    .B(CMD_logic_shift_right),
    .C(_00624_),
    .D(_01229_),
    .X(_01230_));
 sky130_fd_sc_hd__or3_1 _07146_ (.A(_00557_),
    .B(_00631_),
    .C(_01230_),
    .X(_01231_));
 sky130_fd_sc_hd__nand2_1 _07147_ (.A(_01157_),
    .B(CMD_set),
    .Y(_01232_));
 sky130_fd_sc_hd__or4_1 _07148_ (.A(CMD_not),
    .B(_00545_),
    .C(CMD_and),
    .D(_01232_),
    .X(_01233_));
 sky130_fd_sc_hd__or4_1 _07149_ (.A(\shift.left ),
    .B(CMD_logic_shift_right),
    .C(_00624_),
    .D(_01233_),
    .X(_01234_));
 sky130_fd_sc_hd__or4_1 _07150_ (.A(_00557_),
    .B(\current_state[5] ),
    .C(_00634_),
    .D(_01234_),
    .X(_01235_));
 sky130_fd_sc_hd__or4_1 _07151_ (.A(_00528_),
    .B(_00631_),
    .C(_00634_),
    .D(_01171_),
    .X(_01236_));
 sky130_fd_sc_hd__a2111o_1 _07152_ (.A1(_00831_),
    .A2(_00833_),
    .B1(_06264_),
    .C1(_00634_),
    .D1(_01171_),
    .X(_01237_));
 sky130_fd_sc_hd__o2111ai_4 _07153_ (.A1(_00634_),
    .A2(_01231_),
    .B1(_01235_),
    .C1(_01236_),
    .D1(_01237_),
    .Y(_01238_));
 sky130_fd_sc_hd__or2_1 _07154_ (.A(\R2[1] ),
    .B(_01238_),
    .X(_01239_));
 sky130_fd_sc_hd__nand2_1 _07155_ (.A(_01238_),
    .B(_00670_),
    .Y(_01240_));
 sky130_fd_sc_hd__a31o_1 _07156_ (.A1(_01239_),
    .A2(_01214_),
    .A3(_01240_),
    .B1(_01159_),
    .X(_01241_));
 sky130_fd_sc_hd__a2bb2o_1 _07157_ (.A1_N(_01227_),
    .A2_N(_01241_),
    .B1(_00669_),
    .B2(_01159_),
    .X(_01242_));
 sky130_fd_sc_hd__buf_4 _07158_ (.A(_01198_),
    .X(_01243_));
 sky130_fd_sc_hd__inv_2 _07159_ (.A(_01206_),
    .Y(_01244_));
 sky130_fd_sc_hd__buf_4 _07160_ (.A(_01244_),
    .X(_01245_));
 sky130_fd_sc_hd__or4_1 _07161_ (.A(_01159_),
    .B(_01202_),
    .C(_01208_),
    .D(_01190_),
    .X(_01246_));
 sky130_fd_sc_hd__a2111o_1 _07162_ (.A1(_00567_),
    .A2(_01243_),
    .B1(_01220_),
    .C1(_01245_),
    .D1(_01246_),
    .X(_01247_));
 sky130_fd_sc_hd__or2b_2 _07163_ (.A(_01242_),
    .B_N(_01247_),
    .X(_01248_));
 sky130_fd_sc_hd__nor2_4 _07164_ (.A(_01225_),
    .B(_01248_),
    .Y(_01249_));
 sky130_fd_sc_hd__buf_4 _07165_ (.A(_01249_),
    .X(_01250_));
 sky130_fd_sc_hd__mux2_1 _07166_ (.A0(\Oset[3][0] ),
    .A1(_01218_),
    .S(_01250_),
    .X(_01251_));
 sky130_fd_sc_hd__clkbuf_1 _07167_ (.A(_01251_),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _07168_ (.A0(\result_reg_Lshift[1] ),
    .A1(\result_reg_Rshift[1] ),
    .S(_01165_),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _07169_ (.A0(\result_reg_not[1] ),
    .A1(_01252_),
    .S(_01168_),
    .X(_01253_));
 sky130_fd_sc_hd__clkbuf_4 _07170_ (.A(_01190_),
    .X(_01254_));
 sky130_fd_sc_hd__buf_2 _07171_ (.A(_01193_),
    .X(_01255_));
 sky130_fd_sc_hd__or2_1 _07172_ (.A(net8),
    .B(_01255_),
    .X(_01256_));
 sky130_fd_sc_hd__mux2_1 _07173_ (.A0(_00702_),
    .A1(_00703_),
    .S(_01174_),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _07174_ (.A0(_00701_),
    .A1(_01257_),
    .S(_01177_),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _07175_ (.A0(_00700_),
    .A1(_01258_),
    .S(_01182_),
    .X(_01259_));
 sky130_fd_sc_hd__nand2_1 _07176_ (.A(_01259_),
    .B(_01255_),
    .Y(_01260_));
 sky130_fd_sc_hd__nand2_4 _07177_ (.A(_00551_),
    .B(_01243_),
    .Y(_01261_));
 sky130_fd_sc_hd__o21a_1 _07178_ (.A1(\result_reg_and[1] ),
    .A2(_01207_),
    .B1(_01261_),
    .X(_01262_));
 sky130_fd_sc_hd__clkbuf_4 _07179_ (.A(_01204_),
    .X(_01263_));
 sky130_fd_sc_hd__clkbuf_4 _07180_ (.A(_01202_),
    .X(_01264_));
 sky130_fd_sc_hd__inv_2 _07181_ (.A(_01204_),
    .Y(_01265_));
 sky130_fd_sc_hd__clkbuf_4 _07182_ (.A(_01265_),
    .X(_01266_));
 sky130_fd_sc_hd__buf_2 _07183_ (.A(_01264_),
    .X(_01267_));
 sky130_fd_sc_hd__nand2_1 _07184_ (.A(_01267_),
    .B(_00702_),
    .Y(_01268_));
 sky130_fd_sc_hd__o211a_1 _07185_ (.A1(\result_reg_add[1] ),
    .A2(_01264_),
    .B1(_01266_),
    .C1(_01268_),
    .X(_01269_));
 sky130_fd_sc_hd__a211o_1 _07186_ (.A1(\result_reg_mul[1] ),
    .A2(_01263_),
    .B1(_01245_),
    .C1(_01269_),
    .X(_01270_));
 sky130_fd_sc_hd__buf_2 _07187_ (.A(_01261_),
    .X(_01271_));
 sky130_fd_sc_hd__o2bb2a_1 _07188_ (.A1_N(_01262_),
    .A2_N(_01270_),
    .B1(_00708_),
    .B2(_01271_),
    .X(_01272_));
 sky130_fd_sc_hd__o21ai_1 _07189_ (.A1(_01272_),
    .A2(_01238_),
    .B1(_01215_),
    .Y(_01273_));
 sky130_fd_sc_hd__a31o_1 _07190_ (.A1(_01254_),
    .A2(_01256_),
    .A3(_01260_),
    .B1(_01273_),
    .X(_01274_));
 sky130_fd_sc_hd__clkbuf_4 _07191_ (.A(_01220_),
    .X(_01275_));
 sky130_fd_sc_hd__clkbuf_4 _07192_ (.A(_01160_),
    .X(_01276_));
 sky130_fd_sc_hd__a21oi_1 _07193_ (.A1(_00694_),
    .A2(_01275_),
    .B1(_01276_),
    .Y(_01277_));
 sky130_fd_sc_hd__a22o_4 _07194_ (.A1(_01161_),
    .A2(_01253_),
    .B1(_01274_),
    .B2(_01277_),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _07195_ (.A0(\Oset[3][1] ),
    .A1(_01278_),
    .S(_01250_),
    .X(_01279_));
 sky130_fd_sc_hd__clkbuf_1 _07196_ (.A(_01279_),
    .X(_00075_));
 sky130_fd_sc_hd__mux2_1 _07197_ (.A0(\result_reg_Lshift[2] ),
    .A1(\result_reg_Rshift[2] ),
    .S(_01165_),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _07198_ (.A0(\result_reg_not[2] ),
    .A1(_01280_),
    .S(_01168_),
    .X(_01281_));
 sky130_fd_sc_hd__inv_2 _07199_ (.A(\result_reg_and[2] ),
    .Y(_01282_));
 sky130_fd_sc_hd__mux2_1 _07200_ (.A0(\result_reg_add[2] ),
    .A1(\result_reg_sub[2] ),
    .S(_01202_),
    .X(_01283_));
 sky130_fd_sc_hd__nor2_1 _07201_ (.A(_01204_),
    .B(_01283_),
    .Y(_01284_));
 sky130_fd_sc_hd__a211o_1 _07202_ (.A1(_00727_),
    .A2(_01204_),
    .B1(_01245_),
    .C1(_01284_),
    .X(_01285_));
 sky130_fd_sc_hd__o211a_1 _07203_ (.A1(_01282_),
    .A2(_01207_),
    .B1(_01261_),
    .C1(_01285_),
    .X(_01286_));
 sky130_fd_sc_hd__a211o_1 _07204_ (.A1(_00738_),
    .A2(_01208_),
    .B1(_01190_),
    .C1(_01286_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _07205_ (.A0(_00728_),
    .A1(_00729_),
    .S(_01173_),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _07206_ (.A0(_00727_),
    .A1(_01288_),
    .S(_01176_),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _07207_ (.A0(_00726_),
    .A1(_01289_),
    .S(_01181_),
    .X(_01290_));
 sky130_fd_sc_hd__nor2_1 _07208_ (.A(net9),
    .B(_01186_),
    .Y(_01291_));
 sky130_fd_sc_hd__a211o_1 _07209_ (.A1(_01290_),
    .A2(_01193_),
    .B1(_01191_),
    .C1(_01291_),
    .X(_01292_));
 sky130_fd_sc_hd__and3_1 _07210_ (.A(_01287_),
    .B(_01292_),
    .C(_01214_),
    .X(_01293_));
 sky130_fd_sc_hd__a211o_1 _07211_ (.A1(_00724_),
    .A2(_01220_),
    .B1(_01160_),
    .C1(_01293_),
    .X(_01294_));
 sky130_fd_sc_hd__a21bo_4 _07212_ (.A1(_01161_),
    .A2(_01281_),
    .B1_N(_01294_),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _07213_ (.A0(\Oset[3][2] ),
    .A1(_01295_),
    .S(_01250_),
    .X(_01296_));
 sky130_fd_sc_hd__clkbuf_1 _07214_ (.A(_01296_),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _07215_ (.A0(\result_reg_Lshift[3] ),
    .A1(\result_reg_Rshift[3] ),
    .S(_01165_),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _07216_ (.A0(\result_reg_not[3] ),
    .A1(_01297_),
    .S(_01168_),
    .X(_01298_));
 sky130_fd_sc_hd__clkbuf_4 _07217_ (.A(_01207_),
    .X(_01299_));
 sky130_fd_sc_hd__nor2_1 _07218_ (.A(\result_reg_and[3] ),
    .B(_01299_),
    .Y(_01300_));
 sky130_fd_sc_hd__nor2_1 _07219_ (.A(\result_reg_add[3] ),
    .B(_01267_),
    .Y(_01301_));
 sky130_fd_sc_hd__a211o_1 _07220_ (.A1(_00770_),
    .A2(_01267_),
    .B1(_01263_),
    .C1(_01301_),
    .X(_01302_));
 sky130_fd_sc_hd__o211a_1 _07221_ (.A1(_00765_),
    .A2(_01266_),
    .B1(_01299_),
    .C1(_01302_),
    .X(_01303_));
 sky130_fd_sc_hd__o21ai_1 _07222_ (.A1(_01300_),
    .A2(_01303_),
    .B1(_01271_),
    .Y(_01304_));
 sky130_fd_sc_hd__or2_1 _07223_ (.A(\result_reg_or[3] ),
    .B(_01199_),
    .X(_01305_));
 sky130_fd_sc_hd__inv_2 _07224_ (.A(\result_reg_set[3] ),
    .Y(_01306_));
 sky130_fd_sc_hd__mux2_1 _07225_ (.A0(_00770_),
    .A1(_00762_),
    .S(_01174_),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _07226_ (.A0(_00765_),
    .A1(_01307_),
    .S(_01177_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _07227_ (.A0(_01306_),
    .A1(_01308_),
    .S(_01182_),
    .X(_01309_));
 sky130_fd_sc_hd__nand2_1 _07228_ (.A(_01309_),
    .B(_01255_),
    .Y(_01310_));
 sky130_fd_sc_hd__o211a_1 _07229_ (.A1(net10),
    .A2(_01187_),
    .B1(_01254_),
    .C1(_01310_),
    .X(_01311_));
 sky130_fd_sc_hd__a311o_1 _07230_ (.A1(_01192_),
    .A2(_01304_),
    .A3(_01305_),
    .B1(_01275_),
    .C1(_01311_),
    .X(_01312_));
 sky130_fd_sc_hd__a21oi_1 _07231_ (.A1(_00761_),
    .A2(_01275_),
    .B1(_01276_),
    .Y(_01313_));
 sky130_fd_sc_hd__a22o_4 _07232_ (.A1(_01161_),
    .A2(_01298_),
    .B1(_01312_),
    .B2(_01313_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _07233_ (.A0(\Oset[3][3] ),
    .A1(_01314_),
    .S(_01250_),
    .X(_01315_));
 sky130_fd_sc_hd__clkbuf_1 _07234_ (.A(_01315_),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _07235_ (.A0(\result_reg_Lshift[4] ),
    .A1(\result_reg_Rshift[4] ),
    .S(_01165_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _07236_ (.A0(\result_reg_not[4] ),
    .A1(_01316_),
    .S(_01168_),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _07237_ (.A0(_00788_),
    .A1(_00789_),
    .S(_01173_),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _07238_ (.A0(_00787_),
    .A1(_01318_),
    .S(_01176_),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _07239_ (.A0(_00786_),
    .A1(_01319_),
    .S(_01181_),
    .X(_01320_));
 sky130_fd_sc_hd__nor2_1 _07240_ (.A(net11),
    .B(_01193_),
    .Y(_01321_));
 sky130_fd_sc_hd__a211o_1 _07241_ (.A1(_01320_),
    .A2(_01187_),
    .B1(_01192_),
    .C1(_01321_),
    .X(_01322_));
 sky130_fd_sc_hd__inv_2 _07242_ (.A(\result_reg_and[4] ),
    .Y(_01323_));
 sky130_fd_sc_hd__nor2_1 _07243_ (.A(\result_reg_add[4] ),
    .B(_01202_),
    .Y(_01324_));
 sky130_fd_sc_hd__a211o_1 _07244_ (.A1(_00788_),
    .A2(_01202_),
    .B1(_01204_),
    .C1(_01324_),
    .X(_01325_));
 sky130_fd_sc_hd__o211a_1 _07245_ (.A1(_00787_),
    .A2(_01266_),
    .B1(_01207_),
    .C1(_01325_),
    .X(_01326_));
 sky130_fd_sc_hd__a21o_1 _07246_ (.A1(_01323_),
    .A2(_01245_),
    .B1(_01326_),
    .X(_01327_));
 sky130_fd_sc_hd__nor2_1 _07247_ (.A(\result_reg_or[4] ),
    .B(_01199_),
    .Y(_01328_));
 sky130_fd_sc_hd__a211o_1 _07248_ (.A1(_01327_),
    .A2(_01271_),
    .B1(_01254_),
    .C1(_01328_),
    .X(_01329_));
 sky130_fd_sc_hd__nor2_1 _07249_ (.A(\result_reg_mac[4] ),
    .B(_01215_),
    .Y(_01330_));
 sky130_fd_sc_hd__a311o_1 _07250_ (.A1(_01322_),
    .A2(_01215_),
    .A3(_01329_),
    .B1(_01159_),
    .C1(_01330_),
    .X(_01331_));
 sky130_fd_sc_hd__a21bo_4 _07251_ (.A1(_01161_),
    .A2(_01317_),
    .B1_N(_01331_),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _07252_ (.A0(\Oset[3][4] ),
    .A1(_01332_),
    .S(_01250_),
    .X(_01333_));
 sky130_fd_sc_hd__clkbuf_1 _07253_ (.A(_01333_),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _07254_ (.A0(\result_reg_Lshift[5] ),
    .A1(\result_reg_Rshift[5] ),
    .S(_01165_),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _07255_ (.A0(\result_reg_not[5] ),
    .A1(_01334_),
    .S(_01168_),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _07256_ (.A0(_00841_),
    .A1(_00812_),
    .S(_01173_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _07257_ (.A0(_00815_),
    .A1(_01336_),
    .S(_01176_),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _07258_ (.A0(_00840_),
    .A1(_01337_),
    .S(_01181_),
    .X(_01338_));
 sky130_fd_sc_hd__nor2_1 _07259_ (.A(net12),
    .B(_01193_),
    .Y(_01339_));
 sky130_fd_sc_hd__a211o_1 _07260_ (.A1(_01338_),
    .A2(_01187_),
    .B1(_01192_),
    .C1(_01339_),
    .X(_01340_));
 sky130_fd_sc_hd__nand2_1 _07261_ (.A(_01264_),
    .B(_00841_),
    .Y(_01341_));
 sky130_fd_sc_hd__o211a_1 _07262_ (.A1(\result_reg_add[5] ),
    .A2(_01264_),
    .B1(_01265_),
    .C1(_01341_),
    .X(_01342_));
 sky130_fd_sc_hd__a211o_1 _07263_ (.A1(\result_reg_mul[5] ),
    .A2(_01263_),
    .B1(_01245_),
    .C1(_01342_),
    .X(_01343_));
 sky130_fd_sc_hd__o21ai_1 _07264_ (.A1(\result_reg_and[5] ),
    .A2(_01299_),
    .B1(_01343_),
    .Y(_01344_));
 sky130_fd_sc_hd__nor2_1 _07265_ (.A(\result_reg_or[5] ),
    .B(_01199_),
    .Y(_01345_));
 sky130_fd_sc_hd__a211o_1 _07266_ (.A1(_01344_),
    .A2(_01199_),
    .B1(_01190_),
    .C1(_01345_),
    .X(_01346_));
 sky130_fd_sc_hd__nor2_1 _07267_ (.A(\result_reg_mac[5] ),
    .B(_01215_),
    .Y(_01347_));
 sky130_fd_sc_hd__a311o_1 _07268_ (.A1(_01340_),
    .A2(_01214_),
    .A3(_01346_),
    .B1(_01159_),
    .C1(_01347_),
    .X(_01348_));
 sky130_fd_sc_hd__a21bo_4 _07269_ (.A1(_01161_),
    .A2(_01335_),
    .B1_N(_01348_),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_1 _07270_ (.A0(\Oset[3][5] ),
    .A1(_01349_),
    .S(_01250_),
    .X(_01350_));
 sky130_fd_sc_hd__clkbuf_1 _07271_ (.A(_01350_),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _07272_ (.A0(\result_reg_Lshift[6] ),
    .A1(\result_reg_Rshift[6] ),
    .S(_01165_),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _07273_ (.A0(\result_reg_not[6] ),
    .A1(_01351_),
    .S(_01168_),
    .X(_01352_));
 sky130_fd_sc_hd__inv_2 _07274_ (.A(\result_reg_set[6] ),
    .Y(_01353_));
 sky130_fd_sc_hd__mux2_1 _07275_ (.A0(_00865_),
    .A1(_00857_),
    .S(_01173_),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _07276_ (.A0(_00860_),
    .A1(_01354_),
    .S(_01176_),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _07277_ (.A0(_01353_),
    .A1(_01355_),
    .S(_01181_),
    .X(_01356_));
 sky130_fd_sc_hd__nor2_1 _07278_ (.A(net13),
    .B(_01193_),
    .Y(_01357_));
 sky130_fd_sc_hd__a211o_1 _07279_ (.A1(_01356_),
    .A2(_01193_),
    .B1(_01192_),
    .C1(_01357_),
    .X(_01358_));
 sky130_fd_sc_hd__inv_2 _07280_ (.A(\result_reg_and[6] ),
    .Y(_01359_));
 sky130_fd_sc_hd__nor2_1 _07281_ (.A(\result_reg_add[6] ),
    .B(_01202_),
    .Y(_01360_));
 sky130_fd_sc_hd__a211o_1 _07282_ (.A1(_00865_),
    .A2(_01202_),
    .B1(_01204_),
    .C1(_01360_),
    .X(_01361_));
 sky130_fd_sc_hd__o211a_1 _07283_ (.A1(_00860_),
    .A2(_01266_),
    .B1(_01206_),
    .C1(_01361_),
    .X(_01362_));
 sky130_fd_sc_hd__a21o_1 _07284_ (.A1(_01359_),
    .A2(_01245_),
    .B1(_01362_),
    .X(_01363_));
 sky130_fd_sc_hd__nor2_1 _07285_ (.A(\result_reg_or[6] ),
    .B(_01199_),
    .Y(_01364_));
 sky130_fd_sc_hd__a211o_1 _07286_ (.A1(_01363_),
    .A2(_01271_),
    .B1(_01190_),
    .C1(_01364_),
    .X(_01365_));
 sky130_fd_sc_hd__nor2_1 _07287_ (.A(\result_reg_mac[6] ),
    .B(_01215_),
    .Y(_01366_));
 sky130_fd_sc_hd__a311o_1 _07288_ (.A1(_01358_),
    .A2(_01214_),
    .A3(_01365_),
    .B1(_01159_),
    .C1(_01366_),
    .X(_01367_));
 sky130_fd_sc_hd__a21bo_4 _07289_ (.A1(_01161_),
    .A2(_01352_),
    .B1_N(_01367_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _07290_ (.A0(\Oset[3][6] ),
    .A1(_01368_),
    .S(_01250_),
    .X(_01369_));
 sky130_fd_sc_hd__clkbuf_1 _07291_ (.A(_01369_),
    .X(_00080_));
 sky130_fd_sc_hd__mux2_1 _07292_ (.A0(\result_reg_Lshift[7] ),
    .A1(\result_reg_Rshift[7] ),
    .S(_01165_),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _07293_ (.A0(\result_reg_not[7] ),
    .A1(_01370_),
    .S(_01168_),
    .X(_01371_));
 sky130_fd_sc_hd__or2_1 _07294_ (.A(net14),
    .B(_01255_),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_1 _07295_ (.A0(_00883_),
    .A1(_00884_),
    .S(_01174_),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _07296_ (.A0(_00882_),
    .A1(_01373_),
    .S(_01177_),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _07297_ (.A0(_00881_),
    .A1(_01374_),
    .S(_01182_),
    .X(_01375_));
 sky130_fd_sc_hd__nand2_1 _07298_ (.A(_01375_),
    .B(_01255_),
    .Y(_01376_));
 sky130_fd_sc_hd__o21a_1 _07299_ (.A1(\result_reg_and[7] ),
    .A2(_01207_),
    .B1(_01261_),
    .X(_01377_));
 sky130_fd_sc_hd__nand2_1 _07300_ (.A(_01267_),
    .B(_00883_),
    .Y(_01378_));
 sky130_fd_sc_hd__o211a_1 _07301_ (.A1(\result_reg_add[7] ),
    .A2(_01264_),
    .B1(_01266_),
    .C1(_01378_),
    .X(_01379_));
 sky130_fd_sc_hd__a211o_1 _07302_ (.A1(\result_reg_mul[7] ),
    .A2(_01263_),
    .B1(_01245_),
    .C1(_01379_),
    .X(_01380_));
 sky130_fd_sc_hd__o2bb2a_1 _07303_ (.A1_N(_01377_),
    .A2_N(_01380_),
    .B1(_00890_),
    .B2(_01271_),
    .X(_01381_));
 sky130_fd_sc_hd__o21ai_1 _07304_ (.A1(_01381_),
    .A2(_01238_),
    .B1(_01215_),
    .Y(_01382_));
 sky130_fd_sc_hd__a31o_1 _07305_ (.A1(_01254_),
    .A2(_01372_),
    .A3(_01376_),
    .B1(_01382_),
    .X(_01383_));
 sky130_fd_sc_hd__a21oi_1 _07306_ (.A1(_00880_),
    .A2(_01275_),
    .B1(_01276_),
    .Y(_01384_));
 sky130_fd_sc_hd__a22o_4 _07307_ (.A1(_01161_),
    .A2(_01371_),
    .B1(_01383_),
    .B2(_01384_),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _07308_ (.A0(\Oset[3][7] ),
    .A1(_01385_),
    .S(_01250_),
    .X(_01386_));
 sky130_fd_sc_hd__clkbuf_1 _07309_ (.A(_01386_),
    .X(_00081_));
 sky130_fd_sc_hd__mux2_1 _07310_ (.A0(\result_reg_Lshift[8] ),
    .A1(\result_reg_Rshift[8] ),
    .S(_01164_),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _07311_ (.A0(\result_reg_not[8] ),
    .A1(_01387_),
    .S(_01167_),
    .X(_01388_));
 sky130_fd_sc_hd__or2_1 _07312_ (.A(net15),
    .B(_01255_),
    .X(_01389_));
 sky130_fd_sc_hd__inv_2 _07313_ (.A(\result_reg_set[8] ),
    .Y(_01390_));
 sky130_fd_sc_hd__mux2_1 _07314_ (.A0(_00912_),
    .A1(_00906_),
    .S(_01174_),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _07315_ (.A0(_00911_),
    .A1(_01391_),
    .S(_01177_),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_1 _07316_ (.A0(_01390_),
    .A1(_01392_),
    .S(_01182_),
    .X(_01393_));
 sky130_fd_sc_hd__nand2_1 _07317_ (.A(_01393_),
    .B(_01255_),
    .Y(_01394_));
 sky130_fd_sc_hd__mux2_1 _07318_ (.A0(\result_reg_add[8] ),
    .A1(\result_reg_sub[8] ),
    .S(_01264_),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _07319_ (.A0(_01395_),
    .A1(\result_reg_mul[8] ),
    .S(_01263_),
    .X(_01396_));
 sky130_fd_sc_hd__and3_1 _07320_ (.A(_00559_),
    .B(\result_reg_and[8] ),
    .C(_01243_),
    .X(_01397_));
 sky130_fd_sc_hd__a211o_1 _07321_ (.A1(_01396_),
    .A2(_01299_),
    .B1(_01208_),
    .C1(_01397_),
    .X(_01398_));
 sky130_fd_sc_hd__or2_1 _07322_ (.A(\result_reg_or[8] ),
    .B(_01199_),
    .X(_01399_));
 sky130_fd_sc_hd__a31o_1 _07323_ (.A1(_01398_),
    .A2(_01192_),
    .A3(_01399_),
    .B1(_01220_),
    .X(_01400_));
 sky130_fd_sc_hd__a31o_1 _07324_ (.A1(_01254_),
    .A2(_01389_),
    .A3(_01394_),
    .B1(_01400_),
    .X(_01401_));
 sky130_fd_sc_hd__a21oi_1 _07325_ (.A1(_00919_),
    .A2(_01275_),
    .B1(_01276_),
    .Y(_01402_));
 sky130_fd_sc_hd__a22o_4 _07326_ (.A1(_01276_),
    .A2(_01388_),
    .B1(_01401_),
    .B2(_01402_),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _07327_ (.A0(\Oset[3][8] ),
    .A1(_01403_),
    .S(_01250_),
    .X(_01404_));
 sky130_fd_sc_hd__clkbuf_1 _07328_ (.A(_01404_),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _07329_ (.A0(\result_reg_Lshift[9] ),
    .A1(\result_reg_Rshift[9] ),
    .S(_01165_),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _07330_ (.A0(\result_reg_not[9] ),
    .A1(_01405_),
    .S(_01168_),
    .X(_01406_));
 sky130_fd_sc_hd__inv_2 _07331_ (.A(\result_reg_and[9] ),
    .Y(_01407_));
 sky130_fd_sc_hd__mux2_1 _07332_ (.A0(\result_reg_add[9] ),
    .A1(\result_reg_sub[9] ),
    .S(_01201_),
    .X(_01408_));
 sky130_fd_sc_hd__nor2_1 _07333_ (.A(_01204_),
    .B(_01408_),
    .Y(_01409_));
 sky130_fd_sc_hd__a211o_1 _07334_ (.A1(_00931_),
    .A2(_01204_),
    .B1(_01244_),
    .C1(_01409_),
    .X(_01410_));
 sky130_fd_sc_hd__o211a_1 _07335_ (.A1(_01407_),
    .A2(_01207_),
    .B1(_01261_),
    .C1(_01410_),
    .X(_01411_));
 sky130_fd_sc_hd__a211o_1 _07336_ (.A1(_00939_),
    .A2(_01208_),
    .B1(_01190_),
    .C1(_01411_),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _07337_ (.A0(_00932_),
    .A1(_00933_),
    .S(_01173_),
    .X(_01413_));
 sky130_fd_sc_hd__mux2_1 _07338_ (.A0(_00931_),
    .A1(_01413_),
    .S(_01176_),
    .X(_01414_));
 sky130_fd_sc_hd__mux2_1 _07339_ (.A0(_00930_),
    .A1(_01414_),
    .S(_01181_),
    .X(_01415_));
 sky130_fd_sc_hd__nor2_1 _07340_ (.A(net16),
    .B(_01186_),
    .Y(_01416_));
 sky130_fd_sc_hd__a211o_1 _07341_ (.A1(_01415_),
    .A2(_01193_),
    .B1(_01191_),
    .C1(_01416_),
    .X(_01417_));
 sky130_fd_sc_hd__and3_1 _07342_ (.A(_01412_),
    .B(_01417_),
    .C(_01214_),
    .X(_01418_));
 sky130_fd_sc_hd__a211o_1 _07343_ (.A1(_00929_),
    .A2(_01220_),
    .B1(_01160_),
    .C1(_01418_),
    .X(_01419_));
 sky130_fd_sc_hd__a21bo_4 _07344_ (.A1(_01161_),
    .A2(_01406_),
    .B1_N(_01419_),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_1 _07345_ (.A0(\Oset[3][9] ),
    .A1(_01420_),
    .S(_01250_),
    .X(_01421_));
 sky130_fd_sc_hd__clkbuf_1 _07346_ (.A(_01421_),
    .X(_00083_));
 sky130_fd_sc_hd__mux2_1 _07347_ (.A0(\result_reg_Lshift[10] ),
    .A1(\result_reg_Rshift[10] ),
    .S(_01164_),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_1 _07348_ (.A0(\result_reg_not[10] ),
    .A1(_01422_),
    .S(_01167_),
    .X(_01423_));
 sky130_fd_sc_hd__or2_1 _07349_ (.A(net2),
    .B(_01255_),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _07350_ (.A0(_00958_),
    .A1(_00959_),
    .S(_01174_),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_1 _07351_ (.A0(_00957_),
    .A1(_01425_),
    .S(_01177_),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_1 _07352_ (.A0(_00956_),
    .A1(_01426_),
    .S(_01182_),
    .X(_01427_));
 sky130_fd_sc_hd__nand2_1 _07353_ (.A(_01427_),
    .B(_01255_),
    .Y(_01428_));
 sky130_fd_sc_hd__o21a_1 _07354_ (.A1(\result_reg_and[10] ),
    .A2(_01207_),
    .B1(_01261_),
    .X(_01429_));
 sky130_fd_sc_hd__nand2_1 _07355_ (.A(_01264_),
    .B(_00958_),
    .Y(_01430_));
 sky130_fd_sc_hd__o211a_1 _07356_ (.A1(\result_reg_add[10] ),
    .A2(_01264_),
    .B1(_01266_),
    .C1(_01430_),
    .X(_01431_));
 sky130_fd_sc_hd__a211o_1 _07357_ (.A1(\result_reg_mul[10] ),
    .A2(_01263_),
    .B1(_01245_),
    .C1(_01431_),
    .X(_01432_));
 sky130_fd_sc_hd__o2bb2a_1 _07358_ (.A1_N(_01429_),
    .A2_N(_01432_),
    .B1(_00965_),
    .B2(_01271_),
    .X(_01433_));
 sky130_fd_sc_hd__o21ai_1 _07359_ (.A1(_01433_),
    .A2(_01238_),
    .B1(_01215_),
    .Y(_01434_));
 sky130_fd_sc_hd__a31o_1 _07360_ (.A1(_01254_),
    .A2(_01424_),
    .A3(_01428_),
    .B1(_01434_),
    .X(_01435_));
 sky130_fd_sc_hd__a21oi_1 _07361_ (.A1(_00955_),
    .A2(_01275_),
    .B1(_01160_),
    .Y(_01436_));
 sky130_fd_sc_hd__a22o_2 _07362_ (.A1(_01276_),
    .A2(_01423_),
    .B1(_01435_),
    .B2(_01436_),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _07363_ (.A0(\Oset[3][10] ),
    .A1(_01437_),
    .S(_01249_),
    .X(_01438_));
 sky130_fd_sc_hd__clkbuf_1 _07364_ (.A(_01438_),
    .X(_00084_));
 sky130_fd_sc_hd__mux2_1 _07365_ (.A0(\result_reg_Lshift[11] ),
    .A1(\result_reg_Rshift[11] ),
    .S(_01164_),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _07366_ (.A0(\result_reg_not[11] ),
    .A1(_01439_),
    .S(_01167_),
    .X(_01440_));
 sky130_fd_sc_hd__nor2_1 _07367_ (.A(\result_reg_and[11] ),
    .B(_01299_),
    .Y(_01441_));
 sky130_fd_sc_hd__nor2_1 _07368_ (.A(\result_reg_add[11] ),
    .B(_01267_),
    .Y(_01442_));
 sky130_fd_sc_hd__a211o_1 _07369_ (.A1(_00991_),
    .A2(_01267_),
    .B1(_01263_),
    .C1(_01442_),
    .X(_01443_));
 sky130_fd_sc_hd__o211a_1 _07370_ (.A1(_00985_),
    .A2(_01266_),
    .B1(_01299_),
    .C1(_01443_),
    .X(_01444_));
 sky130_fd_sc_hd__o21ai_1 _07371_ (.A1(_01441_),
    .A2(_01444_),
    .B1(_01271_),
    .Y(_01445_));
 sky130_fd_sc_hd__nand2_1 _07372_ (.A(_01208_),
    .B(_00989_),
    .Y(_01446_));
 sky130_fd_sc_hd__inv_2 _07373_ (.A(\result_reg_set[11] ),
    .Y(_01447_));
 sky130_fd_sc_hd__mux2_1 _07374_ (.A0(_00991_),
    .A1(_00982_),
    .S(_01174_),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _07375_ (.A0(_00985_),
    .A1(_01448_),
    .S(_01177_),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _07376_ (.A0(_01447_),
    .A1(_01449_),
    .S(_01182_),
    .X(_01450_));
 sky130_fd_sc_hd__nand2_1 _07377_ (.A(_01450_),
    .B(_01187_),
    .Y(_01451_));
 sky130_fd_sc_hd__o211a_1 _07378_ (.A1(net3),
    .A2(_01187_),
    .B1(_01254_),
    .C1(_01451_),
    .X(_01452_));
 sky130_fd_sc_hd__a311o_1 _07379_ (.A1(_01192_),
    .A2(_01445_),
    .A3(_01446_),
    .B1(_01220_),
    .C1(_01452_),
    .X(_01453_));
 sky130_fd_sc_hd__a21oi_1 _07380_ (.A1(_00981_),
    .A2(_01275_),
    .B1(_01160_),
    .Y(_01454_));
 sky130_fd_sc_hd__a22o_2 _07381_ (.A1(_01276_),
    .A2(_01440_),
    .B1(_01453_),
    .B2(_01454_),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _07382_ (.A0(\Oset[3][11] ),
    .A1(_01455_),
    .S(_01249_),
    .X(_01456_));
 sky130_fd_sc_hd__clkbuf_1 _07383_ (.A(_01456_),
    .X(_00085_));
 sky130_fd_sc_hd__mux2_1 _07384_ (.A0(\result_reg_Lshift[12] ),
    .A1(\result_reg_Rshift[12] ),
    .S(_01164_),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _07385_ (.A0(\result_reg_not[12] ),
    .A1(_01457_),
    .S(_01167_),
    .X(_01458_));
 sky130_fd_sc_hd__nor2_1 _07386_ (.A(\result_reg_and[12] ),
    .B(_01299_),
    .Y(_01459_));
 sky130_fd_sc_hd__nor2_1 _07387_ (.A(\result_reg_add[12] ),
    .B(_01267_),
    .Y(_01460_));
 sky130_fd_sc_hd__a211o_1 _07388_ (.A1(_01016_),
    .A2(_01267_),
    .B1(_01263_),
    .C1(_01460_),
    .X(_01461_));
 sky130_fd_sc_hd__o211a_1 _07389_ (.A1(_01010_),
    .A2(_01266_),
    .B1(_01299_),
    .C1(_01461_),
    .X(_01462_));
 sky130_fd_sc_hd__o21ai_1 _07390_ (.A1(_01459_),
    .A2(_01462_),
    .B1(_01271_),
    .Y(_01463_));
 sky130_fd_sc_hd__nand2_1 _07391_ (.A(_01208_),
    .B(_01014_),
    .Y(_01464_));
 sky130_fd_sc_hd__inv_2 _07392_ (.A(\result_reg_set[12] ),
    .Y(_01465_));
 sky130_fd_sc_hd__mux2_1 _07393_ (.A0(_01016_),
    .A1(_01007_),
    .S(_01174_),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _07394_ (.A0(_01010_),
    .A1(_01466_),
    .S(_01177_),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _07395_ (.A0(_01465_),
    .A1(_01467_),
    .S(_01182_),
    .X(_01468_));
 sky130_fd_sc_hd__nand2_1 _07396_ (.A(_01468_),
    .B(_01187_),
    .Y(_01469_));
 sky130_fd_sc_hd__o211a_1 _07397_ (.A1(net4),
    .A2(_01187_),
    .B1(_01254_),
    .C1(_01469_),
    .X(_01470_));
 sky130_fd_sc_hd__a311o_1 _07398_ (.A1(_01192_),
    .A2(_01463_),
    .A3(_01464_),
    .B1(_01220_),
    .C1(_01470_),
    .X(_01471_));
 sky130_fd_sc_hd__a21oi_1 _07399_ (.A1(_01006_),
    .A2(_01275_),
    .B1(_01160_),
    .Y(_01472_));
 sky130_fd_sc_hd__a22o_2 _07400_ (.A1(_01276_),
    .A2(_01458_),
    .B1(_01471_),
    .B2(_01472_),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _07401_ (.A0(\Oset[3][12] ),
    .A1(_01473_),
    .S(_01249_),
    .X(_01474_));
 sky130_fd_sc_hd__clkbuf_1 _07402_ (.A(_01474_),
    .X(_00086_));
 sky130_fd_sc_hd__mux2_1 _07403_ (.A0(\result_reg_Lshift[13] ),
    .A1(\result_reg_Rshift[13] ),
    .S(_01164_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _07404_ (.A0(\result_reg_not[13] ),
    .A1(_01475_),
    .S(_01167_),
    .X(_01476_));
 sky130_fd_sc_hd__nand2_1 _07405_ (.A(_01185_),
    .B(_01032_),
    .Y(_01477_));
 sky130_fd_sc_hd__mux2_1 _07406_ (.A0(_01035_),
    .A1(_01036_),
    .S(_01174_),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _07407_ (.A0(_01034_),
    .A1(_01478_),
    .S(_01177_),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _07408_ (.A0(_01033_),
    .A1(_01479_),
    .S(_01182_),
    .X(_01480_));
 sky130_fd_sc_hd__nand2_1 _07409_ (.A(_01480_),
    .B(_01255_),
    .Y(_01481_));
 sky130_fd_sc_hd__o21a_1 _07410_ (.A1(\result_reg_and[13] ),
    .A2(_01207_),
    .B1(_01261_),
    .X(_01482_));
 sky130_fd_sc_hd__nand2_1 _07411_ (.A(_01264_),
    .B(_01035_),
    .Y(_01483_));
 sky130_fd_sc_hd__o211a_1 _07412_ (.A1(\result_reg_add[13] ),
    .A2(_01264_),
    .B1(_01266_),
    .C1(_01483_),
    .X(_01484_));
 sky130_fd_sc_hd__a211o_1 _07413_ (.A1(\result_reg_mul[13] ),
    .A2(_01263_),
    .B1(_01245_),
    .C1(_01484_),
    .X(_01485_));
 sky130_fd_sc_hd__o2bb2a_1 _07414_ (.A1_N(_01482_),
    .A2_N(_01485_),
    .B1(_01041_),
    .B2(_01271_),
    .X(_01486_));
 sky130_fd_sc_hd__o21ai_1 _07415_ (.A1(_01486_),
    .A2(_01238_),
    .B1(_01215_),
    .Y(_01487_));
 sky130_fd_sc_hd__a31o_1 _07416_ (.A1(_01254_),
    .A2(_01477_),
    .A3(_01481_),
    .B1(_01487_),
    .X(_01488_));
 sky130_fd_sc_hd__a21oi_1 _07417_ (.A1(_01031_),
    .A2(_01275_),
    .B1(_01160_),
    .Y(_01489_));
 sky130_fd_sc_hd__a22o_2 _07418_ (.A1(_01276_),
    .A2(_01476_),
    .B1(_01488_),
    .B2(_01489_),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _07419_ (.A0(\Oset[3][13] ),
    .A1(_01490_),
    .S(_01249_),
    .X(_01491_));
 sky130_fd_sc_hd__clkbuf_1 _07420_ (.A(_01491_),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _07421_ (.A0(\result_reg_Lshift[14] ),
    .A1(\result_reg_Rshift[14] ),
    .S(_01165_),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _07422_ (.A0(\result_reg_not[14] ),
    .A1(_01492_),
    .S(_01168_),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_1 _07423_ (.A0(_01067_),
    .A1(_01057_),
    .S(_01173_),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _07424_ (.A0(_01060_),
    .A1(_01494_),
    .S(_01176_),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _07425_ (.A0(_01066_),
    .A1(_01495_),
    .S(_01181_),
    .X(_01496_));
 sky130_fd_sc_hd__nor2_1 _07426_ (.A(net6),
    .B(_01193_),
    .Y(_01497_));
 sky130_fd_sc_hd__a211o_1 _07427_ (.A1(_01496_),
    .A2(_01193_),
    .B1(_01191_),
    .C1(_01497_),
    .X(_01498_));
 sky130_fd_sc_hd__inv_2 _07428_ (.A(\result_reg_and[14] ),
    .Y(_01499_));
 sky130_fd_sc_hd__nor2_1 _07429_ (.A(\result_reg_add[14] ),
    .B(_01202_),
    .Y(_01500_));
 sky130_fd_sc_hd__a211o_1 _07430_ (.A1(_01067_),
    .A2(_01202_),
    .B1(_01204_),
    .C1(_01500_),
    .X(_01501_));
 sky130_fd_sc_hd__o211a_1 _07431_ (.A1(_01060_),
    .A2(_01265_),
    .B1(_01206_),
    .C1(_01501_),
    .X(_01502_));
 sky130_fd_sc_hd__a21o_1 _07432_ (.A1(_01499_),
    .A2(_01245_),
    .B1(_01502_),
    .X(_01503_));
 sky130_fd_sc_hd__nor2_1 _07433_ (.A(\result_reg_or[14] ),
    .B(_01199_),
    .Y(_01504_));
 sky130_fd_sc_hd__a211o_1 _07434_ (.A1(_01503_),
    .A2(_01261_),
    .B1(_01190_),
    .C1(_01504_),
    .X(_01505_));
 sky130_fd_sc_hd__nor2_1 _07435_ (.A(\result_reg_mac[14] ),
    .B(_01215_),
    .Y(_01506_));
 sky130_fd_sc_hd__a311o_1 _07436_ (.A1(_01498_),
    .A2(_01214_),
    .A3(_01505_),
    .B1(_01159_),
    .C1(_01506_),
    .X(_01507_));
 sky130_fd_sc_hd__a21bo_1 _07437_ (.A1(_01161_),
    .A2(_01493_),
    .B1_N(_01507_),
    .X(_01508_));
 sky130_fd_sc_hd__mux2_1 _07438_ (.A0(\Oset[3][14] ),
    .A1(_01508_),
    .S(_01249_),
    .X(_01509_));
 sky130_fd_sc_hd__clkbuf_1 _07439_ (.A(_01509_),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _07440_ (.A0(\result_reg_Lshift[15] ),
    .A1(\result_reg_Rshift[15] ),
    .S(_01164_),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _07441_ (.A0(\result_reg_not[15] ),
    .A1(_01510_),
    .S(_01167_),
    .X(_01511_));
 sky130_fd_sc_hd__nor2_1 _07442_ (.A(\result_reg_and[15] ),
    .B(_01299_),
    .Y(_01512_));
 sky130_fd_sc_hd__nor2_1 _07443_ (.A(\result_reg_add[15] ),
    .B(_01267_),
    .Y(_01513_));
 sky130_fd_sc_hd__a211o_1 _07444_ (.A1(_01093_),
    .A2(_01267_),
    .B1(_01263_),
    .C1(_01513_),
    .X(_01514_));
 sky130_fd_sc_hd__o211a_1 _07445_ (.A1(_01086_),
    .A2(_01266_),
    .B1(_01299_),
    .C1(_01514_),
    .X(_01515_));
 sky130_fd_sc_hd__o21ai_1 _07446_ (.A1(_01512_),
    .A2(_01515_),
    .B1(_01271_),
    .Y(_01516_));
 sky130_fd_sc_hd__or2_1 _07447_ (.A(\result_reg_or[15] ),
    .B(_01199_),
    .X(_01517_));
 sky130_fd_sc_hd__mux2_1 _07448_ (.A0(_01093_),
    .A1(_01083_),
    .S(_01174_),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _07449_ (.A0(_01086_),
    .A1(_01518_),
    .S(_01177_),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _07450_ (.A0(_01092_),
    .A1(_01519_),
    .S(_01182_),
    .X(_01520_));
 sky130_fd_sc_hd__nand2_1 _07451_ (.A(_01520_),
    .B(_01187_),
    .Y(_01521_));
 sky130_fd_sc_hd__o211a_1 _07452_ (.A1(net7),
    .A2(_01187_),
    .B1(_01254_),
    .C1(_01521_),
    .X(_01522_));
 sky130_fd_sc_hd__a311o_1 _07453_ (.A1(_01192_),
    .A2(_01516_),
    .A3(_01517_),
    .B1(_01220_),
    .C1(_01522_),
    .X(_01523_));
 sky130_fd_sc_hd__a21oi_1 _07454_ (.A1(_01082_),
    .A2(_01275_),
    .B1(_01160_),
    .Y(_01524_));
 sky130_fd_sc_hd__a22o_1 _07455_ (.A1(_01276_),
    .A2(_01511_),
    .B1(_01523_),
    .B2(_01524_),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _07456_ (.A0(\Oset[3][15] ),
    .A1(_01525_),
    .S(_01249_),
    .X(_01526_));
 sky130_fd_sc_hd__clkbuf_1 _07457_ (.A(_01526_),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _07458_ (.A0(\R2[0] ),
    .A1(net27),
    .S(\current_state[2] ),
    .X(_01527_));
 sky130_fd_sc_hd__and2_1 _07459_ (.A(_01527_),
    .B(_01149_),
    .X(_01528_));
 sky130_fd_sc_hd__clkbuf_1 _07460_ (.A(_01528_),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _07461_ (.A0(\R2[1] ),
    .A1(net28),
    .S(\current_state[2] ),
    .X(_01529_));
 sky130_fd_sc_hd__and2_1 _07462_ (.A(_01529_),
    .B(_01149_),
    .X(_01530_));
 sky130_fd_sc_hd__clkbuf_1 _07463_ (.A(_01530_),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _07464_ (.A0(_00498_),
    .A1(net29),
    .S(\current_state[2] ),
    .X(_01531_));
 sky130_fd_sc_hd__clkbuf_4 _07465_ (.A(_00472_),
    .X(_01532_));
 sky130_fd_sc_hd__and2_1 _07466_ (.A(_01531_),
    .B(_01532_),
    .X(_01533_));
 sky130_fd_sc_hd__clkbuf_1 _07467_ (.A(_01533_),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _07468_ (.A0(\R1[1] ),
    .A1(net30),
    .S(\current_state[2] ),
    .X(_01534_));
 sky130_fd_sc_hd__and2_1 _07469_ (.A(_01534_),
    .B(_01532_),
    .X(_01535_));
 sky130_fd_sc_hd__clkbuf_1 _07470_ (.A(_01535_),
    .X(_00093_));
 sky130_fd_sc_hd__buf_4 _07471_ (.A(Hreg3),
    .X(_01536_));
 sky130_fd_sc_hd__clkbuf_4 _07472_ (.A(_01536_),
    .X(_01537_));
 sky130_fd_sc_hd__buf_4 _07473_ (.A(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__nand2_1 _07474_ (.A(_00472_),
    .B(_01538_),
    .Y(_01539_));
 sky130_fd_sc_hd__nor2_4 _07475_ (.A(_00625_),
    .B(_01539_),
    .Y(_01540_));
 sky130_fd_sc_hd__inv_2 _07476_ (.A(_01540_),
    .Y(_01541_));
 sky130_fd_sc_hd__nand2_1 _07477_ (.A(_00572_),
    .B(Him),
    .Y(_01542_));
 sky130_fd_sc_hd__inv_2 _07478_ (.A(_01542_),
    .Y(_01543_));
 sky130_fd_sc_hd__nand2_4 _07479_ (.A(_00538_),
    .B(_01543_),
    .Y(_01544_));
 sky130_fd_sc_hd__clkbuf_4 _07480_ (.A(_01544_),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _07481_ (.A0(_00610_),
    .A1(_00542_),
    .S(_01545_),
    .X(_01546_));
 sky130_fd_sc_hd__nor2_1 _07482_ (.A(_01542_),
    .B(_00533_),
    .Y(_01547_));
 sky130_fd_sc_hd__inv_2 _07483_ (.A(_01547_),
    .Y(_01548_));
 sky130_fd_sc_hd__buf_2 _07484_ (.A(_01548_),
    .X(_01549_));
 sky130_fd_sc_hd__nand2_1 _07485_ (.A(_01546_),
    .B(_01549_),
    .Y(_01550_));
 sky130_fd_sc_hd__inv_2 _07486_ (.A(_00586_),
    .Y(_01551_));
 sky130_fd_sc_hd__buf_4 _07487_ (.A(_01551_),
    .X(_01552_));
 sky130_fd_sc_hd__clkbuf_4 _07488_ (.A(_01552_),
    .X(_01553_));
 sky130_fd_sc_hd__buf_4 _07489_ (.A(_01553_),
    .X(_01554_));
 sky130_fd_sc_hd__nor2_1 _07490_ (.A(_01554_),
    .B(_00531_),
    .Y(_01555_));
 sky130_fd_sc_hd__inv_2 _07491_ (.A(_01555_),
    .Y(_01556_));
 sky130_fd_sc_hd__nor2_1 _07492_ (.A(_00557_),
    .B(_01556_),
    .Y(_01557_));
 sky130_fd_sc_hd__and2_1 _07493_ (.A(_00550_),
    .B(_00598_),
    .X(_01558_));
 sky130_fd_sc_hd__nand2_2 _07494_ (.A(_01557_),
    .B(_01558_),
    .Y(_01559_));
 sky130_fd_sc_hd__nand2_2 _07495_ (.A(_01557_),
    .B(_01180_),
    .Y(_01560_));
 sky130_fd_sc_hd__buf_2 _07496_ (.A(_01560_),
    .X(_01561_));
 sky130_fd_sc_hd__o211a_1 _07497_ (.A1(\result_reg_mul[0] ),
    .A2(_01549_),
    .B1(_01559_),
    .C1(_01561_),
    .X(_01562_));
 sky130_fd_sc_hd__and3_1 _07498_ (.A(_01557_),
    .B(net1),
    .C(_01558_),
    .X(_01563_));
 sky130_fd_sc_hd__nor2_1 _07499_ (.A(_01170_),
    .B(_01561_),
    .Y(_01564_));
 sky130_fd_sc_hd__a211o_1 _07500_ (.A1(_01550_),
    .A2(_01562_),
    .B1(_01563_),
    .C1(_01564_),
    .X(_01565_));
 sky130_fd_sc_hd__nand2_1 _07501_ (.A(_00569_),
    .B(_01543_),
    .Y(_01566_));
 sky130_fd_sc_hd__and3_1 _07502_ (.A(_01566_),
    .B(_01559_),
    .C(_01560_),
    .X(_01567_));
 sky130_fd_sc_hd__inv_2 _07503_ (.A(_01567_),
    .Y(_01568_));
 sky130_fd_sc_hd__clkbuf_4 _07504_ (.A(_01568_),
    .X(_01569_));
 sky130_fd_sc_hd__clkbuf_4 _07505_ (.A(_01540_),
    .X(_01570_));
 sky130_fd_sc_hd__buf_4 _07506_ (.A(Hreg2),
    .X(_01571_));
 sky130_fd_sc_hd__nand2_4 _07507_ (.A(_01196_),
    .B(_01571_),
    .Y(_01572_));
 sky130_fd_sc_hd__inv_2 _07508_ (.A(_01572_),
    .Y(_01573_));
 sky130_fd_sc_hd__clkbuf_4 _07509_ (.A(_01573_),
    .X(_01574_));
 sky130_fd_sc_hd__nand2_1 _07510_ (.A(_01571_),
    .B(CMD_and),
    .Y(_01575_));
 sky130_fd_sc_hd__or4_1 _07511_ (.A(\shift.left ),
    .B(CMD_logic_shift_right),
    .C(_00624_),
    .D(_01575_),
    .X(_01576_));
 sky130_fd_sc_hd__or4_4 _07512_ (.A(_00557_),
    .B(_00631_),
    .C(_00634_),
    .D(_01576_),
    .X(_01577_));
 sky130_fd_sc_hd__clkinv_4 _07513_ (.A(_01571_),
    .Y(_01578_));
 sky130_fd_sc_hd__nor2_4 _07514_ (.A(_01578_),
    .B(_00537_),
    .Y(_01579_));
 sky130_fd_sc_hd__inv_2 _07515_ (.A(_01579_),
    .Y(_01580_));
 sky130_fd_sc_hd__clkbuf_4 _07516_ (.A(_01580_),
    .X(_01581_));
 sky130_fd_sc_hd__nand2_1 _07517_ (.A(_01581_),
    .B(\result_reg_add[0] ),
    .Y(_01582_));
 sky130_fd_sc_hd__nor2_2 _07518_ (.A(_01578_),
    .B(_00533_),
    .Y(_01583_));
 sky130_fd_sc_hd__inv_2 _07519_ (.A(_01583_),
    .Y(_01584_));
 sky130_fd_sc_hd__clkbuf_4 _07520_ (.A(_01584_),
    .X(_01585_));
 sky130_fd_sc_hd__clkbuf_4 _07521_ (.A(_01579_),
    .X(_01586_));
 sky130_fd_sc_hd__nand2_1 _07522_ (.A(_01586_),
    .B(\result_reg_sub[0] ),
    .Y(_01587_));
 sky130_fd_sc_hd__nand2_1 _07523_ (.A(_00559_),
    .B(_01571_),
    .Y(_01588_));
 sky130_fd_sc_hd__clkbuf_4 _07524_ (.A(_01588_),
    .X(_01589_));
 sky130_fd_sc_hd__o21ai_1 _07525_ (.A1(\result_reg_mul[0] ),
    .A2(_01585_),
    .B1(_01589_),
    .Y(_01590_));
 sky130_fd_sc_hd__a31o_1 _07526_ (.A1(_01582_),
    .A2(_01585_),
    .A3(_01587_),
    .B1(_01590_),
    .X(_01591_));
 sky130_fd_sc_hd__o21ai_1 _07527_ (.A1(_01209_),
    .A2(_01577_),
    .B1(_01591_),
    .Y(_01592_));
 sky130_fd_sc_hd__clkbuf_4 _07528_ (.A(_01567_),
    .X(_01593_));
 sky130_fd_sc_hd__clkbuf_4 _07529_ (.A(_01593_),
    .X(_01594_));
 sky130_fd_sc_hd__clkbuf_4 _07530_ (.A(_01572_),
    .X(_01595_));
 sky130_fd_sc_hd__or2_1 _07531_ (.A(\result_reg_or[0] ),
    .B(_01595_),
    .X(_01596_));
 sky130_fd_sc_hd__o211a_1 _07532_ (.A1(_01574_),
    .A2(_01592_),
    .B1(_01594_),
    .C1(_01596_),
    .X(_01597_));
 sky130_fd_sc_hd__a211o_1 _07533_ (.A1(_01565_),
    .A2(_01569_),
    .B1(_01570_),
    .C1(_01597_),
    .X(_01598_));
 sky130_fd_sc_hd__o21ai_2 _07534_ (.A1(\result_reg_mac[0] ),
    .A2(_01541_),
    .B1(_01598_),
    .Y(_01599_));
 sky130_fd_sc_hd__nor2_4 _07535_ (.A(_00921_),
    .B(_01556_),
    .Y(_01600_));
 sky130_fd_sc_hd__inv_2 _07536_ (.A(_01600_),
    .Y(_01601_));
 sky130_fd_sc_hd__inv_2 _07537_ (.A(_00641_),
    .Y(_01602_));
 sky130_fd_sc_hd__nor2_2 _07538_ (.A(_01602_),
    .B(_01556_),
    .Y(_01603_));
 sky130_fd_sc_hd__inv_2 _07539_ (.A(_01603_),
    .Y(_01604_));
 sky130_fd_sc_hd__nand2_1 _07540_ (.A(_01555_),
    .B(_00640_),
    .Y(_01605_));
 sky130_fd_sc_hd__and3_2 _07541_ (.A(_01601_),
    .B(_01604_),
    .C(_01605_),
    .X(_01606_));
 sky130_fd_sc_hd__clkbuf_4 _07542_ (.A(_01601_),
    .X(_01607_));
 sky130_fd_sc_hd__clkbuf_4 _07543_ (.A(_01603_),
    .X(_01608_));
 sky130_fd_sc_hd__nor2_1 _07544_ (.A(\result_reg_Rshift[0] ),
    .B(_01608_),
    .Y(_01609_));
 sky130_fd_sc_hd__a21o_1 _07545_ (.A1(_01608_),
    .A2(_00659_),
    .B1(_01600_),
    .X(_01610_));
 sky130_fd_sc_hd__inv_2 _07546_ (.A(_01606_),
    .Y(_01611_));
 sky130_fd_sc_hd__buf_4 _07547_ (.A(_01611_),
    .X(_01612_));
 sky130_fd_sc_hd__buf_4 _07548_ (.A(_01612_),
    .X(_01613_));
 sky130_fd_sc_hd__o221a_1 _07549_ (.A1(_00652_),
    .A2(_01607_),
    .B1(_01609_),
    .B2(_01610_),
    .C1(_01613_),
    .X(_01614_));
 sky130_fd_sc_hd__a21oi_4 _07550_ (.A1(_01599_),
    .A2(_01606_),
    .B1(_01614_),
    .Y(_01615_));
 sky130_fd_sc_hd__o21a_1 _07551_ (.A1(\R1[1] ),
    .A2(_01541_),
    .B1(_01606_),
    .X(_01616_));
 sky130_fd_sc_hd__nor2_1 _07552_ (.A(_00670_),
    .B(_01593_),
    .Y(_01617_));
 sky130_fd_sc_hd__a211o_1 _07553_ (.A1(\R2[1] ),
    .A2(_01593_),
    .B1(_01540_),
    .C1(_01617_),
    .X(_01618_));
 sky130_fd_sc_hd__o2bb2a_1 _07554_ (.A1_N(_01616_),
    .A2_N(_01618_),
    .B1(_00669_),
    .B2(_01606_),
    .X(_01619_));
 sky130_fd_sc_hd__or3b_1 _07555_ (.A(_01583_),
    .B(_01573_),
    .C_N(_01588_),
    .X(_01620_));
 sky130_fd_sc_hd__a211o_1 _07556_ (.A1(_01571_),
    .A2(_00565_),
    .B1(_01540_),
    .C1(_01579_),
    .X(_01621_));
 sky130_fd_sc_hd__or4_1 _07557_ (.A(_01611_),
    .B(_01620_),
    .C(_01621_),
    .D(_01568_),
    .X(_01622_));
 sky130_fd_sc_hd__or2b_1 _07558_ (.A(_01619_),
    .B_N(_01622_),
    .X(_01623_));
 sky130_fd_sc_hd__nor2_1 _07559_ (.A(_00681_),
    .B(_01568_),
    .Y(_01624_));
 sky130_fd_sc_hd__a211o_1 _07560_ (.A1(\R0[0] ),
    .A2(_01568_),
    .B1(_01540_),
    .C1(_01624_),
    .X(_01625_));
 sky130_fd_sc_hd__o21a_1 _07561_ (.A1(_00498_),
    .A2(_01541_),
    .B1(_01606_),
    .X(_01626_));
 sky130_fd_sc_hd__a22o_2 _07562_ (.A1(\R3[0] ),
    .A2(_01612_),
    .B1(_01625_),
    .B2(_01626_),
    .X(_01627_));
 sky130_fd_sc_hd__nand2b_4 _07563_ (.A_N(_01623_),
    .B(_01627_),
    .Y(_01628_));
 sky130_fd_sc_hd__clkbuf_8 _07564_ (.A(_01628_),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_1 _07565_ (.A0(_01615_),
    .A1(\H[3][0] ),
    .S(_01629_),
    .X(_01630_));
 sky130_fd_sc_hd__clkbuf_1 _07566_ (.A(_01630_),
    .X(_00094_));
 sky130_fd_sc_hd__nor2_1 _07567_ (.A(_00690_),
    .B(_01608_),
    .Y(_01631_));
 sky130_fd_sc_hd__a211o_1 _07568_ (.A1(\result_reg_Lshift[1] ),
    .A2(_01608_),
    .B1(_01600_),
    .C1(_01631_),
    .X(_01632_));
 sky130_fd_sc_hd__clkbuf_4 _07569_ (.A(_01600_),
    .X(_01633_));
 sky130_fd_sc_hd__nand2_1 _07570_ (.A(_01633_),
    .B(_00689_),
    .Y(_01634_));
 sky130_fd_sc_hd__clkbuf_4 _07571_ (.A(_01559_),
    .X(_01635_));
 sky130_fd_sc_hd__mux2_1 _07572_ (.A0(_00702_),
    .A1(_00703_),
    .S(_01545_),
    .X(_01636_));
 sky130_fd_sc_hd__o21ai_1 _07573_ (.A1(\result_reg_mul[1] ),
    .A2(_01549_),
    .B1(_01561_),
    .Y(_01637_));
 sky130_fd_sc_hd__a21o_1 _07574_ (.A1(_01636_),
    .A2(_01549_),
    .B1(_01637_),
    .X(_01638_));
 sky130_fd_sc_hd__o211ai_1 _07575_ (.A1(_00700_),
    .A2(_01561_),
    .B1(_01635_),
    .C1(_01638_),
    .Y(_01639_));
 sky130_fd_sc_hd__or2_1 _07576_ (.A(net8),
    .B(_01635_),
    .X(_01640_));
 sky130_fd_sc_hd__nand2_1 _07577_ (.A(_01581_),
    .B(\result_reg_add[1] ),
    .Y(_01641_));
 sky130_fd_sc_hd__nand2_1 _07578_ (.A(_01586_),
    .B(\result_reg_sub[1] ),
    .Y(_01642_));
 sky130_fd_sc_hd__o21ai_1 _07579_ (.A1(\result_reg_mul[1] ),
    .A2(_01585_),
    .B1(_01589_),
    .Y(_01643_));
 sky130_fd_sc_hd__a31o_1 _07580_ (.A1(_01641_),
    .A2(_01585_),
    .A3(_01642_),
    .B1(_01643_),
    .X(_01644_));
 sky130_fd_sc_hd__o21ai_1 _07581_ (.A1(_00715_),
    .A2(_01577_),
    .B1(_01644_),
    .Y(_01645_));
 sky130_fd_sc_hd__nand2_1 _07582_ (.A(_01574_),
    .B(_00708_),
    .Y(_01646_));
 sky130_fd_sc_hd__o211a_1 _07583_ (.A1(_01574_),
    .A2(_01645_),
    .B1(_01593_),
    .C1(_01646_),
    .X(_01647_));
 sky130_fd_sc_hd__a311o_1 _07584_ (.A1(_01639_),
    .A2(_01569_),
    .A3(_01640_),
    .B1(_01570_),
    .C1(_01647_),
    .X(_01648_));
 sky130_fd_sc_hd__o21a_1 _07585_ (.A1(\result_reg_mac[1] ),
    .A2(_01541_),
    .B1(_01606_),
    .X(_01649_));
 sky130_fd_sc_hd__a32o_4 _07586_ (.A1(_01613_),
    .A2(_01632_),
    .A3(_01634_),
    .B1(_01648_),
    .B2(_01649_),
    .X(_01650_));
 sky130_fd_sc_hd__mux2_1 _07587_ (.A0(_01650_),
    .A1(\H[3][1] ),
    .S(_01629_),
    .X(_01651_));
 sky130_fd_sc_hd__clkbuf_1 _07588_ (.A(_01651_),
    .X(_00095_));
 sky130_fd_sc_hd__mux2_1 _07589_ (.A0(_00728_),
    .A1(_00729_),
    .S(_01545_),
    .X(_01652_));
 sky130_fd_sc_hd__buf_2 _07590_ (.A(_01548_),
    .X(_01653_));
 sky130_fd_sc_hd__o21ai_1 _07591_ (.A1(\result_reg_mul[2] ),
    .A2(_01653_),
    .B1(_01561_),
    .Y(_01654_));
 sky130_fd_sc_hd__a21o_1 _07592_ (.A1(_01652_),
    .A2(_01549_),
    .B1(_01654_),
    .X(_01655_));
 sky130_fd_sc_hd__buf_2 _07593_ (.A(_01560_),
    .X(_01656_));
 sky130_fd_sc_hd__or2_1 _07594_ (.A(_00726_),
    .B(_01656_),
    .X(_01657_));
 sky130_fd_sc_hd__clkbuf_4 _07595_ (.A(_01559_),
    .X(_01658_));
 sky130_fd_sc_hd__nor2_1 _07596_ (.A(net9),
    .B(_01658_),
    .Y(_01659_));
 sky130_fd_sc_hd__a31o_1 _07597_ (.A1(_01655_),
    .A2(_01635_),
    .A3(_01657_),
    .B1(_01659_),
    .X(_01660_));
 sky130_fd_sc_hd__nand2_1 _07598_ (.A(_01581_),
    .B(\result_reg_add[2] ),
    .Y(_01661_));
 sky130_fd_sc_hd__nand2_1 _07599_ (.A(_01586_),
    .B(\result_reg_sub[2] ),
    .Y(_01662_));
 sky130_fd_sc_hd__clkbuf_4 _07600_ (.A(_01584_),
    .X(_01663_));
 sky130_fd_sc_hd__o21ai_1 _07601_ (.A1(\result_reg_mul[2] ),
    .A2(_01663_),
    .B1(_01589_),
    .Y(_01664_));
 sky130_fd_sc_hd__a31o_1 _07602_ (.A1(_01661_),
    .A2(_01585_),
    .A3(_01662_),
    .B1(_01664_),
    .X(_01665_));
 sky130_fd_sc_hd__clkbuf_4 _07603_ (.A(_01571_),
    .X(_01666_));
 sky130_fd_sc_hd__clkbuf_4 _07604_ (.A(_01588_),
    .X(_01667_));
 sky130_fd_sc_hd__o2bb2a_1 _07605_ (.A1_N(_01666_),
    .A2_N(_00551_),
    .B1(_01282_),
    .B2(_01667_),
    .X(_01668_));
 sky130_fd_sc_hd__a221o_1 _07606_ (.A1(_00738_),
    .A2(_01574_),
    .B1(_01665_),
    .B2(_01668_),
    .C1(_01569_),
    .X(_01669_));
 sky130_fd_sc_hd__o21ai_1 _07607_ (.A1(_01594_),
    .A2(_01660_),
    .B1(_01669_),
    .Y(_01670_));
 sky130_fd_sc_hd__mux2_1 _07608_ (.A0(_01670_),
    .A1(\result_reg_mac[2] ),
    .S(_01570_),
    .X(_01671_));
 sky130_fd_sc_hd__clkbuf_4 _07609_ (.A(_01603_),
    .X(_01672_));
 sky130_fd_sc_hd__nand2_1 _07610_ (.A(_01608_),
    .B(_00755_),
    .Y(_01673_));
 sky130_fd_sc_hd__o211a_1 _07611_ (.A1(\result_reg_Rshift[2] ),
    .A2(_01672_),
    .B1(_01607_),
    .C1(_01673_),
    .X(_01674_));
 sky130_fd_sc_hd__a21o_1 _07612_ (.A1(\result_reg_not[2] ),
    .A2(_01633_),
    .B1(_01674_),
    .X(_01675_));
 sky130_fd_sc_hd__mux2_4 _07613_ (.A0(_01671_),
    .A1(_01675_),
    .S(_01613_),
    .X(_01676_));
 sky130_fd_sc_hd__mux2_1 _07614_ (.A0(_01676_),
    .A1(\H[3][2] ),
    .S(_01629_),
    .X(_01677_));
 sky130_fd_sc_hd__clkbuf_1 _07615_ (.A(_01677_),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_1 _07616_ (.A0(_00770_),
    .A1(_00762_),
    .S(_01545_),
    .X(_01678_));
 sky130_fd_sc_hd__clkbuf_4 _07617_ (.A(_01548_),
    .X(_01679_));
 sky130_fd_sc_hd__o21ai_1 _07618_ (.A1(\result_reg_mul[3] ),
    .A2(_01679_),
    .B1(_01561_),
    .Y(_01680_));
 sky130_fd_sc_hd__a21o_1 _07619_ (.A1(_01678_),
    .A2(_01549_),
    .B1(_01680_),
    .X(_01681_));
 sky130_fd_sc_hd__buf_2 _07620_ (.A(_01560_),
    .X(_01682_));
 sky130_fd_sc_hd__or2_1 _07621_ (.A(_01306_),
    .B(_01682_),
    .X(_01683_));
 sky130_fd_sc_hd__nor2_1 _07622_ (.A(net10),
    .B(_01658_),
    .Y(_01684_));
 sky130_fd_sc_hd__a31o_1 _07623_ (.A1(_01681_),
    .A2(_01635_),
    .A3(_01683_),
    .B1(_01684_),
    .X(_01685_));
 sky130_fd_sc_hd__nand2_1 _07624_ (.A(_01581_),
    .B(\result_reg_add[3] ),
    .Y(_01686_));
 sky130_fd_sc_hd__nand2_1 _07625_ (.A(_01586_),
    .B(\result_reg_sub[3] ),
    .Y(_01687_));
 sky130_fd_sc_hd__clkbuf_4 _07626_ (.A(_01584_),
    .X(_01688_));
 sky130_fd_sc_hd__o21ai_1 _07627_ (.A1(\result_reg_mul[3] ),
    .A2(_01688_),
    .B1(_01667_),
    .Y(_01689_));
 sky130_fd_sc_hd__a31o_1 _07628_ (.A1(_01686_),
    .A2(_01663_),
    .A3(_01687_),
    .B1(_01689_),
    .X(_01690_));
 sky130_fd_sc_hd__inv_2 _07629_ (.A(_01577_),
    .Y(_01691_));
 sky130_fd_sc_hd__nand2_1 _07630_ (.A(_01691_),
    .B(\result_reg_and[3] ),
    .Y(_01692_));
 sky130_fd_sc_hd__nor2_1 _07631_ (.A(\result_reg_or[3] ),
    .B(_01595_),
    .Y(_01693_));
 sky130_fd_sc_hd__a311o_1 _07632_ (.A1(_01690_),
    .A2(_01595_),
    .A3(_01692_),
    .B1(_01569_),
    .C1(_01693_),
    .X(_01694_));
 sky130_fd_sc_hd__o21ai_1 _07633_ (.A1(_01594_),
    .A2(_01685_),
    .B1(_01694_),
    .Y(_01695_));
 sky130_fd_sc_hd__mux2_1 _07634_ (.A0(_01695_),
    .A1(\result_reg_mac[3] ),
    .S(_01570_),
    .X(_01696_));
 sky130_fd_sc_hd__nand2_1 _07635_ (.A(_01608_),
    .B(_00779_),
    .Y(_01697_));
 sky130_fd_sc_hd__o211a_1 _07636_ (.A1(\result_reg_Rshift[3] ),
    .A2(_01672_),
    .B1(_01607_),
    .C1(_01697_),
    .X(_01698_));
 sky130_fd_sc_hd__a21o_1 _07637_ (.A1(\result_reg_not[3] ),
    .A2(_01633_),
    .B1(_01698_),
    .X(_01699_));
 sky130_fd_sc_hd__mux2_4 _07638_ (.A0(_01696_),
    .A1(_01699_),
    .S(_01613_),
    .X(_01700_));
 sky130_fd_sc_hd__mux2_1 _07639_ (.A0(_01700_),
    .A1(\H[3][3] ),
    .S(_01629_),
    .X(_01701_));
 sky130_fd_sc_hd__clkbuf_1 _07640_ (.A(_01701_),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _07641_ (.A0(_00788_),
    .A1(_00789_),
    .S(_01545_),
    .X(_01702_));
 sky130_fd_sc_hd__o21ai_1 _07642_ (.A1(\result_reg_mul[4] ),
    .A2(_01679_),
    .B1(_01561_),
    .Y(_01703_));
 sky130_fd_sc_hd__a21o_1 _07643_ (.A1(_01702_),
    .A2(_01549_),
    .B1(_01703_),
    .X(_01704_));
 sky130_fd_sc_hd__or2_1 _07644_ (.A(_00786_),
    .B(_01682_),
    .X(_01705_));
 sky130_fd_sc_hd__nor2_1 _07645_ (.A(net11),
    .B(_01658_),
    .Y(_01706_));
 sky130_fd_sc_hd__a31o_1 _07646_ (.A1(_01704_),
    .A2(_01635_),
    .A3(_01705_),
    .B1(_01706_),
    .X(_01707_));
 sky130_fd_sc_hd__nand2_1 _07647_ (.A(_01581_),
    .B(\result_reg_add[4] ),
    .Y(_01708_));
 sky130_fd_sc_hd__nand2_1 _07648_ (.A(_01586_),
    .B(\result_reg_sub[4] ),
    .Y(_01709_));
 sky130_fd_sc_hd__o21ai_1 _07649_ (.A1(\result_reg_mul[4] ),
    .A2(_01688_),
    .B1(_01589_),
    .Y(_01710_));
 sky130_fd_sc_hd__a31o_1 _07650_ (.A1(_01708_),
    .A2(_01585_),
    .A3(_01709_),
    .B1(_01710_),
    .X(_01711_));
 sky130_fd_sc_hd__o2bb2a_1 _07651_ (.A1_N(_01571_),
    .A2_N(_00551_),
    .B1(_01323_),
    .B2(_01667_),
    .X(_01712_));
 sky130_fd_sc_hd__a221o_1 _07652_ (.A1(_00795_),
    .A2(_01574_),
    .B1(_01711_),
    .B2(_01712_),
    .C1(_01569_),
    .X(_01713_));
 sky130_fd_sc_hd__o21ai_1 _07653_ (.A1(_01594_),
    .A2(_01707_),
    .B1(_01713_),
    .Y(_01714_));
 sky130_fd_sc_hd__mux2_1 _07654_ (.A0(_01714_),
    .A1(\result_reg_mac[4] ),
    .S(_01570_),
    .X(_01715_));
 sky130_fd_sc_hd__clkbuf_4 _07655_ (.A(_01603_),
    .X(_01716_));
 sky130_fd_sc_hd__nand2_1 _07656_ (.A(_01716_),
    .B(_00806_),
    .Y(_01717_));
 sky130_fd_sc_hd__o211a_1 _07657_ (.A1(\result_reg_Rshift[4] ),
    .A2(_01672_),
    .B1(_01607_),
    .C1(_01717_),
    .X(_01718_));
 sky130_fd_sc_hd__a21o_1 _07658_ (.A1(\result_reg_not[4] ),
    .A2(_01633_),
    .B1(_01718_),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_4 _07659_ (.A0(_01715_),
    .A1(_01719_),
    .S(_01613_),
    .X(_01720_));
 sky130_fd_sc_hd__mux2_1 _07660_ (.A0(_01720_),
    .A1(\H[3][4] ),
    .S(_01629_),
    .X(_01721_));
 sky130_fd_sc_hd__clkbuf_1 _07661_ (.A(_01721_),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _07662_ (.A0(_00841_),
    .A1(_00812_),
    .S(_01545_),
    .X(_01722_));
 sky130_fd_sc_hd__o21ai_1 _07663_ (.A1(\result_reg_mul[5] ),
    .A2(_01679_),
    .B1(_01561_),
    .Y(_01723_));
 sky130_fd_sc_hd__a21o_1 _07664_ (.A1(_01722_),
    .A2(_01549_),
    .B1(_01723_),
    .X(_01724_));
 sky130_fd_sc_hd__or2_1 _07665_ (.A(_00840_),
    .B(_01682_),
    .X(_01725_));
 sky130_fd_sc_hd__nor2_1 _07666_ (.A(net12),
    .B(_01658_),
    .Y(_01726_));
 sky130_fd_sc_hd__a31o_1 _07667_ (.A1(_01724_),
    .A2(_01635_),
    .A3(_01725_),
    .B1(_01726_),
    .X(_01727_));
 sky130_fd_sc_hd__nand2_1 _07668_ (.A(_01580_),
    .B(\result_reg_add[5] ),
    .Y(_01728_));
 sky130_fd_sc_hd__nand2_1 _07669_ (.A(_01579_),
    .B(\result_reg_sub[5] ),
    .Y(_01729_));
 sky130_fd_sc_hd__o21ai_1 _07670_ (.A1(\result_reg_mul[5] ),
    .A2(_01688_),
    .B1(_01667_),
    .Y(_01730_));
 sky130_fd_sc_hd__a31o_1 _07671_ (.A1(_01728_),
    .A2(_01663_),
    .A3(_01729_),
    .B1(_01730_),
    .X(_01731_));
 sky130_fd_sc_hd__nand2_1 _07672_ (.A(_01691_),
    .B(\result_reg_and[5] ),
    .Y(_01732_));
 sky130_fd_sc_hd__nor2_1 _07673_ (.A(\result_reg_or[5] ),
    .B(_01595_),
    .Y(_01733_));
 sky130_fd_sc_hd__a311o_1 _07674_ (.A1(_01731_),
    .A2(_01572_),
    .A3(_01732_),
    .B1(_01568_),
    .C1(_01733_),
    .X(_01734_));
 sky130_fd_sc_hd__o21ai_1 _07675_ (.A1(_01594_),
    .A2(_01727_),
    .B1(_01734_),
    .Y(_01735_));
 sky130_fd_sc_hd__mux2_1 _07676_ (.A0(_01735_),
    .A1(\result_reg_mac[5] ),
    .S(_01570_),
    .X(_01736_));
 sky130_fd_sc_hd__nand2_1 _07677_ (.A(_01716_),
    .B(_00850_),
    .Y(_01737_));
 sky130_fd_sc_hd__o211a_1 _07678_ (.A1(\result_reg_Rshift[5] ),
    .A2(_01672_),
    .B1(_01607_),
    .C1(_01737_),
    .X(_01738_));
 sky130_fd_sc_hd__a21o_1 _07679_ (.A1(\result_reg_not[5] ),
    .A2(_01633_),
    .B1(_01738_),
    .X(_01739_));
 sky130_fd_sc_hd__mux2_4 _07680_ (.A0(_01736_),
    .A1(_01739_),
    .S(_01613_),
    .X(_01740_));
 sky130_fd_sc_hd__mux2_1 _07681_ (.A0(_01740_),
    .A1(\H[3][5] ),
    .S(_01629_),
    .X(_01741_));
 sky130_fd_sc_hd__clkbuf_1 _07682_ (.A(_01741_),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _07683_ (.A0(_00865_),
    .A1(_00857_),
    .S(_01545_),
    .X(_01742_));
 sky130_fd_sc_hd__o21ai_1 _07684_ (.A1(\result_reg_mul[6] ),
    .A2(_01679_),
    .B1(_01656_),
    .Y(_01743_));
 sky130_fd_sc_hd__a21o_1 _07685_ (.A1(_01742_),
    .A2(_01549_),
    .B1(_01743_),
    .X(_01744_));
 sky130_fd_sc_hd__or2_1 _07686_ (.A(_01353_),
    .B(_01682_),
    .X(_01745_));
 sky130_fd_sc_hd__clkbuf_4 _07687_ (.A(_01559_),
    .X(_01746_));
 sky130_fd_sc_hd__nor2_1 _07688_ (.A(net13),
    .B(_01746_),
    .Y(_01747_));
 sky130_fd_sc_hd__a31o_1 _07689_ (.A1(_01744_),
    .A2(_01635_),
    .A3(_01745_),
    .B1(_01747_),
    .X(_01748_));
 sky130_fd_sc_hd__nand2_1 _07690_ (.A(_01580_),
    .B(\result_reg_add[6] ),
    .Y(_01749_));
 sky130_fd_sc_hd__nand2_1 _07691_ (.A(_01579_),
    .B(\result_reg_sub[6] ),
    .Y(_01750_));
 sky130_fd_sc_hd__o21ai_1 _07692_ (.A1(\result_reg_mul[6] ),
    .A2(_01688_),
    .B1(_01667_),
    .Y(_01751_));
 sky130_fd_sc_hd__a31o_1 _07693_ (.A1(_01749_),
    .A2(_01663_),
    .A3(_01750_),
    .B1(_01751_),
    .X(_01752_));
 sky130_fd_sc_hd__nand2_1 _07694_ (.A(_01691_),
    .B(\result_reg_and[6] ),
    .Y(_01753_));
 sky130_fd_sc_hd__nor2_1 _07695_ (.A(\result_reg_or[6] ),
    .B(_01595_),
    .Y(_01754_));
 sky130_fd_sc_hd__a311o_1 _07696_ (.A1(_01752_),
    .A2(_01572_),
    .A3(_01753_),
    .B1(_01568_),
    .C1(_01754_),
    .X(_01755_));
 sky130_fd_sc_hd__o21ai_1 _07697_ (.A1(_01594_),
    .A2(_01748_),
    .B1(_01755_),
    .Y(_01756_));
 sky130_fd_sc_hd__mux2_1 _07698_ (.A0(_01756_),
    .A1(\result_reg_mac[6] ),
    .S(_01570_),
    .X(_01757_));
 sky130_fd_sc_hd__nand2_1 _07699_ (.A(_01716_),
    .B(_00874_),
    .Y(_01758_));
 sky130_fd_sc_hd__o211a_1 _07700_ (.A1(\result_reg_Rshift[6] ),
    .A2(_01672_),
    .B1(_01607_),
    .C1(_01758_),
    .X(_01759_));
 sky130_fd_sc_hd__a21o_1 _07701_ (.A1(\result_reg_not[6] ),
    .A2(_01633_),
    .B1(_01759_),
    .X(_01760_));
 sky130_fd_sc_hd__mux2_4 _07702_ (.A0(_01757_),
    .A1(_01760_),
    .S(_01613_),
    .X(_01761_));
 sky130_fd_sc_hd__mux2_1 _07703_ (.A0(_01761_),
    .A1(\H[3][6] ),
    .S(_01629_),
    .X(_01762_));
 sky130_fd_sc_hd__clkbuf_1 _07704_ (.A(_01762_),
    .X(_00100_));
 sky130_fd_sc_hd__nor2_1 _07705_ (.A(\result_reg_Rshift[7] ),
    .B(_01608_),
    .Y(_01763_));
 sky130_fd_sc_hd__a211o_1 _07706_ (.A1(_00901_),
    .A2(_01608_),
    .B1(_01600_),
    .C1(_01763_),
    .X(_01764_));
 sky130_fd_sc_hd__o21ai_1 _07707_ (.A1(_00899_),
    .A2(_01607_),
    .B1(_01764_),
    .Y(_01765_));
 sky130_fd_sc_hd__mux2_1 _07708_ (.A0(_00883_),
    .A1(_00884_),
    .S(_01545_),
    .X(_01766_));
 sky130_fd_sc_hd__o21ai_1 _07709_ (.A1(\result_reg_mul[7] ),
    .A2(_01653_),
    .B1(_01561_),
    .Y(_01767_));
 sky130_fd_sc_hd__a21o_1 _07710_ (.A1(_01766_),
    .A2(_01549_),
    .B1(_01767_),
    .X(_01768_));
 sky130_fd_sc_hd__or2_1 _07711_ (.A(_00881_),
    .B(_01561_),
    .X(_01769_));
 sky130_fd_sc_hd__nor2_1 _07712_ (.A(net14),
    .B(_01635_),
    .Y(_01770_));
 sky130_fd_sc_hd__a311o_1 _07713_ (.A1(_01768_),
    .A2(_01635_),
    .A3(_01769_),
    .B1(_01593_),
    .C1(_01770_),
    .X(_01771_));
 sky130_fd_sc_hd__nand2_1 _07714_ (.A(_01581_),
    .B(\result_reg_add[7] ),
    .Y(_01772_));
 sky130_fd_sc_hd__nand2_1 _07715_ (.A(_01586_),
    .B(\result_reg_sub[7] ),
    .Y(_01773_));
 sky130_fd_sc_hd__o21ai_1 _07716_ (.A1(\result_reg_mul[7] ),
    .A2(_01585_),
    .B1(_01589_),
    .Y(_01774_));
 sky130_fd_sc_hd__a31o_1 _07717_ (.A1(_01772_),
    .A2(_01585_),
    .A3(_01773_),
    .B1(_01774_),
    .X(_01775_));
 sky130_fd_sc_hd__inv_2 _07718_ (.A(\result_reg_and[7] ),
    .Y(_01776_));
 sky130_fd_sc_hd__o2bb2a_1 _07719_ (.A1_N(_01666_),
    .A2_N(_00551_),
    .B1(_01776_),
    .B2(_01589_),
    .X(_01777_));
 sky130_fd_sc_hd__a221o_1 _07720_ (.A1(_00890_),
    .A2(_01574_),
    .B1(_01775_),
    .B2(_01777_),
    .C1(_01569_),
    .X(_01778_));
 sky130_fd_sc_hd__a31o_1 _07721_ (.A1(_01771_),
    .A2(_01541_),
    .A3(_01778_),
    .B1(_01612_),
    .X(_01779_));
 sky130_fd_sc_hd__a21oi_1 _07722_ (.A1(_00880_),
    .A2(_01570_),
    .B1(_01779_),
    .Y(_01780_));
 sky130_fd_sc_hd__a21o_2 _07723_ (.A1(_01613_),
    .A2(_01765_),
    .B1(_01780_),
    .X(_01781_));
 sky130_fd_sc_hd__mux2_1 _07724_ (.A0(_01781_),
    .A1(\H[3][7] ),
    .S(_01629_),
    .X(_01782_));
 sky130_fd_sc_hd__clkbuf_1 _07725_ (.A(_01782_),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _07726_ (.A0(_00912_),
    .A1(_00906_),
    .S(_01545_),
    .X(_01783_));
 sky130_fd_sc_hd__o21ai_1 _07727_ (.A1(\result_reg_mul[8] ),
    .A2(_01679_),
    .B1(_01656_),
    .Y(_01784_));
 sky130_fd_sc_hd__a21o_1 _07728_ (.A1(_01783_),
    .A2(_01653_),
    .B1(_01784_),
    .X(_01785_));
 sky130_fd_sc_hd__or2_1 _07729_ (.A(_01390_),
    .B(_01682_),
    .X(_01786_));
 sky130_fd_sc_hd__nor2_1 _07730_ (.A(net15),
    .B(_01746_),
    .Y(_01787_));
 sky130_fd_sc_hd__a31o_1 _07731_ (.A1(_01785_),
    .A2(_01635_),
    .A3(_01786_),
    .B1(_01787_),
    .X(_01788_));
 sky130_fd_sc_hd__nand2_1 _07732_ (.A(_01580_),
    .B(\result_reg_add[8] ),
    .Y(_01789_));
 sky130_fd_sc_hd__nand2_1 _07733_ (.A(_01579_),
    .B(\result_reg_sub[8] ),
    .Y(_01790_));
 sky130_fd_sc_hd__o21ai_1 _07734_ (.A1(\result_reg_mul[8] ),
    .A2(_01688_),
    .B1(_01667_),
    .Y(_01791_));
 sky130_fd_sc_hd__a31o_1 _07735_ (.A1(_01789_),
    .A2(_01663_),
    .A3(_01790_),
    .B1(_01791_),
    .X(_01792_));
 sky130_fd_sc_hd__nand2_1 _07736_ (.A(_01691_),
    .B(\result_reg_and[8] ),
    .Y(_01793_));
 sky130_fd_sc_hd__nor2_1 _07737_ (.A(\result_reg_or[8] ),
    .B(_01595_),
    .Y(_01794_));
 sky130_fd_sc_hd__a311o_1 _07738_ (.A1(_01792_),
    .A2(_01572_),
    .A3(_01793_),
    .B1(_01568_),
    .C1(_01794_),
    .X(_01795_));
 sky130_fd_sc_hd__o21ai_1 _07739_ (.A1(_01594_),
    .A2(_01788_),
    .B1(_01795_),
    .Y(_01796_));
 sky130_fd_sc_hd__mux2_1 _07740_ (.A0(_01796_),
    .A1(\result_reg_mac[8] ),
    .S(_01570_),
    .X(_01797_));
 sky130_fd_sc_hd__nand2_1 _07741_ (.A(_01716_),
    .B(_00923_),
    .Y(_01798_));
 sky130_fd_sc_hd__o211a_1 _07742_ (.A1(\result_reg_Rshift[8] ),
    .A2(_01672_),
    .B1(_01607_),
    .C1(_01798_),
    .X(_01799_));
 sky130_fd_sc_hd__a21o_1 _07743_ (.A1(\result_reg_not[8] ),
    .A2(_01633_),
    .B1(_01799_),
    .X(_01800_));
 sky130_fd_sc_hd__mux2_2 _07744_ (.A0(_01797_),
    .A1(_01800_),
    .S(_01613_),
    .X(_01801_));
 sky130_fd_sc_hd__mux2_1 _07745_ (.A0(_01801_),
    .A1(\H[3][8] ),
    .S(_01629_),
    .X(_01802_));
 sky130_fd_sc_hd__clkbuf_1 _07746_ (.A(_01802_),
    .X(_00102_));
 sky130_fd_sc_hd__nor2_1 _07747_ (.A(\result_reg_mac[9] ),
    .B(_01541_),
    .Y(_01803_));
 sky130_fd_sc_hd__mux2_1 _07748_ (.A0(\result_reg_add[9] ),
    .A1(\result_reg_sub[9] ),
    .S(_01579_),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_1 _07749_ (.A0(_01804_),
    .A1(\result_reg_mul[9] ),
    .S(_01583_),
    .X(_01805_));
 sky130_fd_sc_hd__nand2_1 _07750_ (.A(_01805_),
    .B(_01589_),
    .Y(_01806_));
 sky130_fd_sc_hd__o211a_1 _07751_ (.A1(_01407_),
    .A2(_01577_),
    .B1(_01572_),
    .C1(_01806_),
    .X(_01807_));
 sky130_fd_sc_hd__a211o_1 _07752_ (.A1(_00939_),
    .A2(_01574_),
    .B1(_01569_),
    .C1(_01807_),
    .X(_01808_));
 sky130_fd_sc_hd__mux2_1 _07753_ (.A0(_00932_),
    .A1(_00933_),
    .S(_01544_),
    .X(_01809_));
 sky130_fd_sc_hd__o21ai_1 _07754_ (.A1(\result_reg_mul[9] ),
    .A2(_01548_),
    .B1(_01656_),
    .Y(_01810_));
 sky130_fd_sc_hd__a21o_1 _07755_ (.A1(_01809_),
    .A2(_01653_),
    .B1(_01810_),
    .X(_01811_));
 sky130_fd_sc_hd__or2_1 _07756_ (.A(_00930_),
    .B(_01560_),
    .X(_01812_));
 sky130_fd_sc_hd__nor2_1 _07757_ (.A(net16),
    .B(_01746_),
    .Y(_01813_));
 sky130_fd_sc_hd__a311o_1 _07758_ (.A1(_01811_),
    .A2(_01746_),
    .A3(_01812_),
    .B1(_01593_),
    .C1(_01813_),
    .X(_01814_));
 sky130_fd_sc_hd__a31o_1 _07759_ (.A1(_01808_),
    .A2(_01541_),
    .A3(_01814_),
    .B1(_01612_),
    .X(_01815_));
 sky130_fd_sc_hd__nor2_1 _07760_ (.A(\result_reg_Rshift[9] ),
    .B(_01608_),
    .Y(_01816_));
 sky130_fd_sc_hd__a211o_1 _07761_ (.A1(_00949_),
    .A2(_01608_),
    .B1(_01600_),
    .C1(_01816_),
    .X(_01817_));
 sky130_fd_sc_hd__o21ai_1 _07762_ (.A1(_00948_),
    .A2(_01607_),
    .B1(_01817_),
    .Y(_01818_));
 sky130_fd_sc_hd__a2bb2o_2 _07763_ (.A1_N(_01803_),
    .A2_N(_01815_),
    .B1(_01613_),
    .B2(_01818_),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_1 _07764_ (.A0(_01819_),
    .A1(\H[3][9] ),
    .S(_01629_),
    .X(_01820_));
 sky130_fd_sc_hd__clkbuf_1 _07765_ (.A(_01820_),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _07766_ (.A0(_00958_),
    .A1(_00959_),
    .S(_01545_),
    .X(_01821_));
 sky130_fd_sc_hd__o21ai_1 _07767_ (.A1(\result_reg_mul[10] ),
    .A2(_01679_),
    .B1(_01656_),
    .Y(_01822_));
 sky130_fd_sc_hd__a21o_1 _07768_ (.A1(_01821_),
    .A2(_01653_),
    .B1(_01822_),
    .X(_01823_));
 sky130_fd_sc_hd__or2_1 _07769_ (.A(_00956_),
    .B(_01682_),
    .X(_01824_));
 sky130_fd_sc_hd__nor2_1 _07770_ (.A(net2),
    .B(_01746_),
    .Y(_01825_));
 sky130_fd_sc_hd__a31o_1 _07771_ (.A1(_01823_),
    .A2(_01658_),
    .A3(_01824_),
    .B1(_01825_),
    .X(_01826_));
 sky130_fd_sc_hd__nand2_1 _07772_ (.A(_01581_),
    .B(\result_reg_add[10] ),
    .Y(_01827_));
 sky130_fd_sc_hd__nand2_1 _07773_ (.A(_01586_),
    .B(\result_reg_sub[10] ),
    .Y(_01828_));
 sky130_fd_sc_hd__o21ai_1 _07774_ (.A1(\result_reg_mul[10] ),
    .A2(_01688_),
    .B1(_01589_),
    .Y(_01829_));
 sky130_fd_sc_hd__a31o_1 _07775_ (.A1(_01827_),
    .A2(_01663_),
    .A3(_01828_),
    .B1(_01829_),
    .X(_01830_));
 sky130_fd_sc_hd__inv_2 _07776_ (.A(\result_reg_and[10] ),
    .Y(_01831_));
 sky130_fd_sc_hd__o2bb2a_1 _07777_ (.A1_N(_01571_),
    .A2_N(_00551_),
    .B1(_01831_),
    .B2(_01667_),
    .X(_01832_));
 sky130_fd_sc_hd__a221o_1 _07778_ (.A1(_00965_),
    .A2(_01574_),
    .B1(_01830_),
    .B2(_01832_),
    .C1(_01569_),
    .X(_01833_));
 sky130_fd_sc_hd__o21ai_1 _07779_ (.A1(_01594_),
    .A2(_01826_),
    .B1(_01833_),
    .Y(_01834_));
 sky130_fd_sc_hd__mux2_1 _07780_ (.A0(_01834_),
    .A1(\result_reg_mac[10] ),
    .S(_01570_),
    .X(_01835_));
 sky130_fd_sc_hd__nand2_1 _07781_ (.A(_01716_),
    .B(_00975_),
    .Y(_01836_));
 sky130_fd_sc_hd__o211a_1 _07782_ (.A1(\result_reg_Rshift[10] ),
    .A2(_01672_),
    .B1(_01607_),
    .C1(_01836_),
    .X(_01837_));
 sky130_fd_sc_hd__a21o_1 _07783_ (.A1(\result_reg_not[10] ),
    .A2(_01633_),
    .B1(_01837_),
    .X(_01838_));
 sky130_fd_sc_hd__mux2_2 _07784_ (.A0(_01835_),
    .A1(_01838_),
    .S(_01612_),
    .X(_01839_));
 sky130_fd_sc_hd__mux2_1 _07785_ (.A0(_01839_),
    .A1(\H[3][10] ),
    .S(_01628_),
    .X(_01840_));
 sky130_fd_sc_hd__clkbuf_1 _07786_ (.A(_01840_),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _07787_ (.A0(_00991_),
    .A1(_00982_),
    .S(_01544_),
    .X(_01841_));
 sky130_fd_sc_hd__o21ai_1 _07788_ (.A1(\result_reg_mul[11] ),
    .A2(_01679_),
    .B1(_01656_),
    .Y(_01842_));
 sky130_fd_sc_hd__a21o_1 _07789_ (.A1(_01841_),
    .A2(_01653_),
    .B1(_01842_),
    .X(_01843_));
 sky130_fd_sc_hd__or2_1 _07790_ (.A(_01447_),
    .B(_01682_),
    .X(_01844_));
 sky130_fd_sc_hd__nor2_1 _07791_ (.A(net3),
    .B(_01746_),
    .Y(_01845_));
 sky130_fd_sc_hd__a31o_1 _07792_ (.A1(_01843_),
    .A2(_01658_),
    .A3(_01844_),
    .B1(_01845_),
    .X(_01846_));
 sky130_fd_sc_hd__nand2_1 _07793_ (.A(_01581_),
    .B(\result_reg_add[11] ),
    .Y(_01847_));
 sky130_fd_sc_hd__nand2_1 _07794_ (.A(_01586_),
    .B(\result_reg_sub[11] ),
    .Y(_01848_));
 sky130_fd_sc_hd__o21ai_1 _07795_ (.A1(\result_reg_mul[11] ),
    .A2(_01688_),
    .B1(_01589_),
    .Y(_01849_));
 sky130_fd_sc_hd__a31o_1 _07796_ (.A1(_01847_),
    .A2(_01663_),
    .A3(_01848_),
    .B1(_01849_),
    .X(_01850_));
 sky130_fd_sc_hd__inv_2 _07797_ (.A(\result_reg_and[11] ),
    .Y(_01851_));
 sky130_fd_sc_hd__o2bb2a_1 _07798_ (.A1_N(_01571_),
    .A2_N(_00551_),
    .B1(_01851_),
    .B2(_01588_),
    .X(_01852_));
 sky130_fd_sc_hd__a221o_1 _07799_ (.A1(_00989_),
    .A2(_01574_),
    .B1(_01850_),
    .B2(_01852_),
    .C1(_01569_),
    .X(_01853_));
 sky130_fd_sc_hd__o21ai_1 _07800_ (.A1(_01594_),
    .A2(_01846_),
    .B1(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__mux2_1 _07801_ (.A0(_01854_),
    .A1(\result_reg_mac[11] ),
    .S(_01540_),
    .X(_01855_));
 sky130_fd_sc_hd__nand2_1 _07802_ (.A(_01716_),
    .B(_01000_),
    .Y(_01856_));
 sky130_fd_sc_hd__o211a_1 _07803_ (.A1(\result_reg_Rshift[11] ),
    .A2(_01672_),
    .B1(_01601_),
    .C1(_01856_),
    .X(_01857_));
 sky130_fd_sc_hd__a21o_1 _07804_ (.A1(\result_reg_not[11] ),
    .A2(_01633_),
    .B1(_01857_),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_2 _07805_ (.A0(_01855_),
    .A1(_01858_),
    .S(_01612_),
    .X(_01859_));
 sky130_fd_sc_hd__mux2_1 _07806_ (.A0(_01859_),
    .A1(\H[3][11] ),
    .S(_01628_),
    .X(_01860_));
 sky130_fd_sc_hd__clkbuf_1 _07807_ (.A(_01860_),
    .X(_00105_));
 sky130_fd_sc_hd__mux2_1 _07808_ (.A0(_01016_),
    .A1(_01007_),
    .S(_01544_),
    .X(_01861_));
 sky130_fd_sc_hd__o21ai_1 _07809_ (.A1(\result_reg_mul[12] ),
    .A2(_01679_),
    .B1(_01656_),
    .Y(_01862_));
 sky130_fd_sc_hd__a21o_1 _07810_ (.A1(_01861_),
    .A2(_01653_),
    .B1(_01862_),
    .X(_01863_));
 sky130_fd_sc_hd__or2_1 _07811_ (.A(_01465_),
    .B(_01682_),
    .X(_01864_));
 sky130_fd_sc_hd__nor2_1 _07812_ (.A(net4),
    .B(_01746_),
    .Y(_01865_));
 sky130_fd_sc_hd__a31o_1 _07813_ (.A1(_01863_),
    .A2(_01658_),
    .A3(_01864_),
    .B1(_01865_),
    .X(_01866_));
 sky130_fd_sc_hd__nand2_1 _07814_ (.A(_01581_),
    .B(\result_reg_add[12] ),
    .Y(_01867_));
 sky130_fd_sc_hd__nand2_1 _07815_ (.A(_01586_),
    .B(\result_reg_sub[12] ),
    .Y(_01868_));
 sky130_fd_sc_hd__o21ai_1 _07816_ (.A1(\result_reg_mul[12] ),
    .A2(_01585_),
    .B1(_01589_),
    .Y(_01869_));
 sky130_fd_sc_hd__a31o_1 _07817_ (.A1(_01867_),
    .A2(_01585_),
    .A3(_01868_),
    .B1(_01869_),
    .X(_01870_));
 sky130_fd_sc_hd__nand2_1 _07818_ (.A(_01691_),
    .B(\result_reg_and[12] ),
    .Y(_01871_));
 sky130_fd_sc_hd__o21ai_1 _07819_ (.A1(\result_reg_or[12] ),
    .A2(_01595_),
    .B1(_01593_),
    .Y(_01872_));
 sky130_fd_sc_hd__a31o_1 _07820_ (.A1(_01870_),
    .A2(_01595_),
    .A3(_01871_),
    .B1(_01872_),
    .X(_01873_));
 sky130_fd_sc_hd__o21ai_1 _07821_ (.A1(_01594_),
    .A2(_01866_),
    .B1(_01873_),
    .Y(_01874_));
 sky130_fd_sc_hd__mux2_1 _07822_ (.A0(_01874_),
    .A1(\result_reg_mac[12] ),
    .S(_01540_),
    .X(_01875_));
 sky130_fd_sc_hd__nand2_1 _07823_ (.A(_01716_),
    .B(_01025_),
    .Y(_01876_));
 sky130_fd_sc_hd__o211a_1 _07824_ (.A1(\result_reg_Rshift[12] ),
    .A2(_01672_),
    .B1(_01601_),
    .C1(_01876_),
    .X(_01877_));
 sky130_fd_sc_hd__a21o_1 _07825_ (.A1(\result_reg_not[12] ),
    .A2(_01633_),
    .B1(_01877_),
    .X(_01878_));
 sky130_fd_sc_hd__mux2_1 _07826_ (.A0(_01875_),
    .A1(_01878_),
    .S(_01612_),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_1 _07827_ (.A0(_01879_),
    .A1(\H[3][12] ),
    .S(_01628_),
    .X(_01880_));
 sky130_fd_sc_hd__clkbuf_1 _07828_ (.A(_01880_),
    .X(_00106_));
 sky130_fd_sc_hd__mux2_1 _07829_ (.A0(_01035_),
    .A1(_01036_),
    .S(_01544_),
    .X(_01881_));
 sky130_fd_sc_hd__o21ai_1 _07830_ (.A1(\result_reg_mul[13] ),
    .A2(_01679_),
    .B1(_01656_),
    .Y(_01882_));
 sky130_fd_sc_hd__a21o_1 _07831_ (.A1(_01881_),
    .A2(_01653_),
    .B1(_01882_),
    .X(_01883_));
 sky130_fd_sc_hd__or2_1 _07832_ (.A(_01033_),
    .B(_01682_),
    .X(_01884_));
 sky130_fd_sc_hd__nor2_1 _07833_ (.A(net5),
    .B(_01746_),
    .Y(_01885_));
 sky130_fd_sc_hd__a31o_1 _07834_ (.A1(_01883_),
    .A2(_01658_),
    .A3(_01884_),
    .B1(_01885_),
    .X(_01886_));
 sky130_fd_sc_hd__nand2_1 _07835_ (.A(_01581_),
    .B(\result_reg_add[13] ),
    .Y(_01887_));
 sky130_fd_sc_hd__nand2_1 _07836_ (.A(_01586_),
    .B(\result_reg_sub[13] ),
    .Y(_01888_));
 sky130_fd_sc_hd__o21ai_1 _07837_ (.A1(\result_reg_mul[13] ),
    .A2(_01688_),
    .B1(_01667_),
    .Y(_01889_));
 sky130_fd_sc_hd__a31o_1 _07838_ (.A1(_01887_),
    .A2(_01663_),
    .A3(_01888_),
    .B1(_01889_),
    .X(_01890_));
 sky130_fd_sc_hd__o2bb2a_1 _07839_ (.A1_N(_01571_),
    .A2_N(_00551_),
    .B1(_01042_),
    .B2(_01588_),
    .X(_01891_));
 sky130_fd_sc_hd__a221o_1 _07840_ (.A1(_01041_),
    .A2(_01574_),
    .B1(_01890_),
    .B2(_01891_),
    .C1(_01569_),
    .X(_01892_));
 sky130_fd_sc_hd__o21ai_1 _07841_ (.A1(_01593_),
    .A2(_01886_),
    .B1(_01892_),
    .Y(_01893_));
 sky130_fd_sc_hd__mux2_1 _07842_ (.A0(_01893_),
    .A1(\result_reg_mac[13] ),
    .S(_01540_),
    .X(_01894_));
 sky130_fd_sc_hd__nand2_1 _07843_ (.A(_01716_),
    .B(_01050_),
    .Y(_01895_));
 sky130_fd_sc_hd__o211a_1 _07844_ (.A1(\result_reg_Rshift[13] ),
    .A2(_01672_),
    .B1(_01601_),
    .C1(_01895_),
    .X(_01896_));
 sky130_fd_sc_hd__a21o_1 _07845_ (.A1(\result_reg_not[13] ),
    .A2(_01600_),
    .B1(_01896_),
    .X(_01897_));
 sky130_fd_sc_hd__mux2_1 _07846_ (.A0(_01894_),
    .A1(_01897_),
    .S(_01612_),
    .X(_01898_));
 sky130_fd_sc_hd__mux2_1 _07847_ (.A0(_01898_),
    .A1(\H[3][13] ),
    .S(_01628_),
    .X(_01899_));
 sky130_fd_sc_hd__clkbuf_1 _07848_ (.A(_01899_),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _07849_ (.A0(_01067_),
    .A1(_01057_),
    .S(_01544_),
    .X(_01900_));
 sky130_fd_sc_hd__o21ai_1 _07850_ (.A1(\result_reg_mul[14] ),
    .A2(_01679_),
    .B1(_01656_),
    .Y(_01901_));
 sky130_fd_sc_hd__a21o_1 _07851_ (.A1(_01900_),
    .A2(_01653_),
    .B1(_01901_),
    .X(_01902_));
 sky130_fd_sc_hd__or2_1 _07852_ (.A(_01066_),
    .B(_01682_),
    .X(_01903_));
 sky130_fd_sc_hd__nor2_1 _07853_ (.A(net6),
    .B(_01746_),
    .Y(_01904_));
 sky130_fd_sc_hd__a31o_1 _07854_ (.A1(_01902_),
    .A2(_01658_),
    .A3(_01903_),
    .B1(_01904_),
    .X(_01905_));
 sky130_fd_sc_hd__nand2_1 _07855_ (.A(_01580_),
    .B(\result_reg_add[14] ),
    .Y(_01906_));
 sky130_fd_sc_hd__nand2_1 _07856_ (.A(_01579_),
    .B(\result_reg_sub[14] ),
    .Y(_01907_));
 sky130_fd_sc_hd__o21ai_1 _07857_ (.A1(\result_reg_mul[14] ),
    .A2(_01688_),
    .B1(_01667_),
    .Y(_01908_));
 sky130_fd_sc_hd__a31o_1 _07858_ (.A1(_01906_),
    .A2(_01663_),
    .A3(_01907_),
    .B1(_01908_),
    .X(_01909_));
 sky130_fd_sc_hd__nand2_1 _07859_ (.A(_01691_),
    .B(\result_reg_and[14] ),
    .Y(_01910_));
 sky130_fd_sc_hd__nor2_1 _07860_ (.A(\result_reg_or[14] ),
    .B(_01595_),
    .Y(_01911_));
 sky130_fd_sc_hd__a311o_1 _07861_ (.A1(_01909_),
    .A2(_01572_),
    .A3(_01910_),
    .B1(_01568_),
    .C1(_01911_),
    .X(_01912_));
 sky130_fd_sc_hd__o21ai_1 _07862_ (.A1(_01593_),
    .A2(_01905_),
    .B1(_01912_),
    .Y(_01913_));
 sky130_fd_sc_hd__mux2_1 _07863_ (.A0(_01913_),
    .A1(\result_reg_mac[14] ),
    .S(_01540_),
    .X(_01914_));
 sky130_fd_sc_hd__nand2_1 _07864_ (.A(_01716_),
    .B(_01076_),
    .Y(_01915_));
 sky130_fd_sc_hd__o211a_1 _07865_ (.A1(\result_reg_Rshift[14] ),
    .A2(_01603_),
    .B1(_01601_),
    .C1(_01915_),
    .X(_01916_));
 sky130_fd_sc_hd__a21o_1 _07866_ (.A1(\result_reg_not[14] ),
    .A2(_01600_),
    .B1(_01916_),
    .X(_01917_));
 sky130_fd_sc_hd__mux2_1 _07867_ (.A0(_01914_),
    .A1(_01917_),
    .S(_01612_),
    .X(_01918_));
 sky130_fd_sc_hd__mux2_1 _07868_ (.A0(_01918_),
    .A1(\H[3][14] ),
    .S(_01628_),
    .X(_01919_));
 sky130_fd_sc_hd__clkbuf_1 _07869_ (.A(_01919_),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _07870_ (.A0(_01093_),
    .A1(_01083_),
    .S(_01544_),
    .X(_01920_));
 sky130_fd_sc_hd__o21ai_1 _07871_ (.A1(\result_reg_mul[15] ),
    .A2(_01548_),
    .B1(_01656_),
    .Y(_01921_));
 sky130_fd_sc_hd__a21o_1 _07872_ (.A1(_01920_),
    .A2(_01653_),
    .B1(_01921_),
    .X(_01922_));
 sky130_fd_sc_hd__or2_1 _07873_ (.A(_01092_),
    .B(_01560_),
    .X(_01923_));
 sky130_fd_sc_hd__nor2_1 _07874_ (.A(net7),
    .B(_01746_),
    .Y(_01924_));
 sky130_fd_sc_hd__a31o_1 _07875_ (.A1(_01922_),
    .A2(_01658_),
    .A3(_01923_),
    .B1(_01924_),
    .X(_01925_));
 sky130_fd_sc_hd__nand2_1 _07876_ (.A(_01580_),
    .B(\result_reg_add[15] ),
    .Y(_01926_));
 sky130_fd_sc_hd__nand2_1 _07877_ (.A(_01579_),
    .B(\result_reg_sub[15] ),
    .Y(_01927_));
 sky130_fd_sc_hd__o21ai_1 _07878_ (.A1(\result_reg_mul[15] ),
    .A2(_01688_),
    .B1(_01667_),
    .Y(_01928_));
 sky130_fd_sc_hd__a31o_1 _07879_ (.A1(_01926_),
    .A2(_01663_),
    .A3(_01927_),
    .B1(_01928_),
    .X(_01929_));
 sky130_fd_sc_hd__nand2_1 _07880_ (.A(_01691_),
    .B(\result_reg_and[15] ),
    .Y(_01930_));
 sky130_fd_sc_hd__nor2_1 _07881_ (.A(\result_reg_or[15] ),
    .B(_01595_),
    .Y(_01931_));
 sky130_fd_sc_hd__a311o_1 _07882_ (.A1(_01929_),
    .A2(_01572_),
    .A3(_01930_),
    .B1(_01568_),
    .C1(_01931_),
    .X(_01932_));
 sky130_fd_sc_hd__o21ai_1 _07883_ (.A1(_01593_),
    .A2(_01925_),
    .B1(_01932_),
    .Y(_01933_));
 sky130_fd_sc_hd__mux2_1 _07884_ (.A0(_01933_),
    .A1(\result_reg_mac[15] ),
    .S(_01540_),
    .X(_01934_));
 sky130_fd_sc_hd__nand2_1 _07885_ (.A(_01716_),
    .B(_01103_),
    .Y(_01935_));
 sky130_fd_sc_hd__o211a_1 _07886_ (.A1(\result_reg_Rshift[15] ),
    .A2(_01603_),
    .B1(_01601_),
    .C1(_01935_),
    .X(_01936_));
 sky130_fd_sc_hd__a21o_1 _07887_ (.A1(\result_reg_not[15] ),
    .A2(_01600_),
    .B1(_01936_),
    .X(_01937_));
 sky130_fd_sc_hd__mux2_1 _07888_ (.A0(_01934_),
    .A1(_01937_),
    .S(_01612_),
    .X(_01938_));
 sky130_fd_sc_hd__mux2_1 _07889_ (.A0(_01938_),
    .A1(\H[3][15] ),
    .S(_01628_),
    .X(_01939_));
 sky130_fd_sc_hd__clkbuf_1 _07890_ (.A(_01939_),
    .X(_00109_));
 sky130_fd_sc_hd__inv_2 _07891_ (.A(_01225_),
    .Y(_01940_));
 sky130_fd_sc_hd__nor2_4 _07892_ (.A(_01940_),
    .B(_01248_),
    .Y(_01941_));
 sky130_fd_sc_hd__buf_4 _07893_ (.A(_01941_),
    .X(_01942_));
 sky130_fd_sc_hd__mux2_1 _07894_ (.A0(\Oset[2][0] ),
    .A1(_01218_),
    .S(_01942_),
    .X(_01943_));
 sky130_fd_sc_hd__clkbuf_1 _07895_ (.A(_01943_),
    .X(_00110_));
 sky130_fd_sc_hd__mux2_1 _07896_ (.A0(\Oset[2][1] ),
    .A1(_01278_),
    .S(_01942_),
    .X(_01944_));
 sky130_fd_sc_hd__clkbuf_1 _07897_ (.A(_01944_),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_1 _07898_ (.A0(\Oset[2][2] ),
    .A1(_01295_),
    .S(_01942_),
    .X(_01945_));
 sky130_fd_sc_hd__clkbuf_1 _07899_ (.A(_01945_),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_1 _07900_ (.A0(\Oset[2][3] ),
    .A1(_01314_),
    .S(_01942_),
    .X(_01946_));
 sky130_fd_sc_hd__clkbuf_1 _07901_ (.A(_01946_),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _07902_ (.A0(\Oset[2][4] ),
    .A1(_01332_),
    .S(_01942_),
    .X(_01947_));
 sky130_fd_sc_hd__clkbuf_1 _07903_ (.A(_01947_),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_1 _07904_ (.A0(\Oset[2][5] ),
    .A1(_01349_),
    .S(_01942_),
    .X(_01948_));
 sky130_fd_sc_hd__clkbuf_1 _07905_ (.A(_01948_),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_1 _07906_ (.A0(\Oset[2][6] ),
    .A1(_01368_),
    .S(_01942_),
    .X(_01949_));
 sky130_fd_sc_hd__clkbuf_1 _07907_ (.A(_01949_),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _07908_ (.A0(\Oset[2][7] ),
    .A1(_01385_),
    .S(_01942_),
    .X(_01950_));
 sky130_fd_sc_hd__clkbuf_1 _07909_ (.A(_01950_),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_1 _07910_ (.A0(\Oset[2][8] ),
    .A1(_01403_),
    .S(_01942_),
    .X(_01951_));
 sky130_fd_sc_hd__clkbuf_1 _07911_ (.A(_01951_),
    .X(_00118_));
 sky130_fd_sc_hd__mux2_1 _07912_ (.A0(\Oset[2][9] ),
    .A1(_01420_),
    .S(_01942_),
    .X(_01952_));
 sky130_fd_sc_hd__clkbuf_1 _07913_ (.A(_01952_),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _07914_ (.A0(\Oset[2][10] ),
    .A1(_01437_),
    .S(_01941_),
    .X(_01953_));
 sky130_fd_sc_hd__clkbuf_1 _07915_ (.A(_01953_),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _07916_ (.A0(\Oset[2][11] ),
    .A1(_01455_),
    .S(_01941_),
    .X(_01954_));
 sky130_fd_sc_hd__clkbuf_1 _07917_ (.A(_01954_),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _07918_ (.A0(\Oset[2][12] ),
    .A1(_01473_),
    .S(_01941_),
    .X(_01955_));
 sky130_fd_sc_hd__clkbuf_1 _07919_ (.A(_01955_),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_1 _07920_ (.A0(\Oset[2][13] ),
    .A1(_01490_),
    .S(_01941_),
    .X(_01956_));
 sky130_fd_sc_hd__clkbuf_1 _07921_ (.A(_01956_),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_1 _07922_ (.A0(\Oset[2][14] ),
    .A1(_01508_),
    .S(_01941_),
    .X(_01957_));
 sky130_fd_sc_hd__clkbuf_1 _07923_ (.A(_01957_),
    .X(_00124_));
 sky130_fd_sc_hd__mux2_1 _07924_ (.A0(\Oset[2][15] ),
    .A1(_01525_),
    .S(_01941_),
    .X(_01958_));
 sky130_fd_sc_hd__clkbuf_1 _07925_ (.A(_01958_),
    .X(_00125_));
 sky130_fd_sc_hd__inv_2 _07926_ (.A(\R3[0] ),
    .Y(_01959_));
 sky130_fd_sc_hd__clkbuf_4 _07927_ (.A(CMD_setloop),
    .X(_01960_));
 sky130_fd_sc_hd__mux2_1 _07928_ (.A0(\LC[0] ),
    .A1(_01959_),
    .S(_01960_),
    .X(_01961_));
 sky130_fd_sc_hd__inv_2 _07929_ (.A(CMD_setloop),
    .Y(_01962_));
 sky130_fd_sc_hd__nand2_1 _07930_ (.A(_06284_),
    .B(_01962_),
    .Y(_01963_));
 sky130_fd_sc_hd__nand2_4 _07931_ (.A(_01963_),
    .B(_00474_),
    .Y(_01964_));
 sky130_fd_sc_hd__nand2_1 _07932_ (.A(_01964_),
    .B(\LC[0] ),
    .Y(_01965_));
 sky130_fd_sc_hd__o21ai_1 _07933_ (.A1(_01961_),
    .A2(_01964_),
    .B1(_01965_),
    .Y(_00126_));
 sky130_fd_sc_hd__nand2_1 _07934_ (.A(\LC[1] ),
    .B(\LC[0] ),
    .Y(_01966_));
 sky130_fd_sc_hd__nand2_1 _07935_ (.A(_06273_),
    .B(_01966_),
    .Y(_01967_));
 sky130_fd_sc_hd__mux2_1 _07936_ (.A0(_01967_),
    .A1(\R3[1] ),
    .S(_01960_),
    .X(_01968_));
 sky130_fd_sc_hd__mux2_1 _07937_ (.A0(_01968_),
    .A1(\LC[1] ),
    .S(_01964_),
    .X(_01969_));
 sky130_fd_sc_hd__clkbuf_1 _07938_ (.A(_01969_),
    .X(_00127_));
 sky130_fd_sc_hd__nand2_1 _07939_ (.A(_06273_),
    .B(\LC[2] ),
    .Y(_01970_));
 sky130_fd_sc_hd__nand2_1 _07940_ (.A(_06274_),
    .B(_01970_),
    .Y(_01971_));
 sky130_fd_sc_hd__mux2_1 _07941_ (.A0(_01971_),
    .A1(\R2[0] ),
    .S(_01960_),
    .X(_01972_));
 sky130_fd_sc_hd__mux2_1 _07942_ (.A0(_01972_),
    .A1(\LC[2] ),
    .S(_01964_),
    .X(_01973_));
 sky130_fd_sc_hd__clkbuf_1 _07943_ (.A(_01973_),
    .X(_00128_));
 sky130_fd_sc_hd__nand2_1 _07944_ (.A(_06274_),
    .B(\LC[3] ),
    .Y(_01974_));
 sky130_fd_sc_hd__and3_1 _07945_ (.A(_06275_),
    .B(_01962_),
    .C(_01974_),
    .X(_01975_));
 sky130_fd_sc_hd__a21oi_1 _07946_ (.A1(_01960_),
    .A2(_00671_),
    .B1(_01975_),
    .Y(_01976_));
 sky130_fd_sc_hd__mux2_1 _07947_ (.A0(_01976_),
    .A1(\LC[3] ),
    .S(_01964_),
    .X(_01977_));
 sky130_fd_sc_hd__clkbuf_1 _07948_ (.A(_01977_),
    .X(_00129_));
 sky130_fd_sc_hd__and2_1 _07949_ (.A(_06275_),
    .B(\LC[4] ),
    .X(_01978_));
 sky130_fd_sc_hd__nand2_1 _07950_ (.A(_06277_),
    .B(_01962_),
    .Y(_01979_));
 sky130_fd_sc_hd__o22a_1 _07951_ (.A1(_00498_),
    .A2(_01962_),
    .B1(_01978_),
    .B2(_01979_),
    .X(_01980_));
 sky130_fd_sc_hd__mux2_1 _07952_ (.A0(_01980_),
    .A1(\LC[4] ),
    .S(_01964_),
    .X(_01981_));
 sky130_fd_sc_hd__clkbuf_1 _07953_ (.A(_01981_),
    .X(_00130_));
 sky130_fd_sc_hd__nand2_1 _07954_ (.A(_06277_),
    .B(\LC[5] ),
    .Y(_01982_));
 sky130_fd_sc_hd__a21o_1 _07955_ (.A1(_06279_),
    .A2(_01982_),
    .B1(_01960_),
    .X(_01983_));
 sky130_fd_sc_hd__o21ai_1 _07956_ (.A1(_01962_),
    .A2(_01226_),
    .B1(_01983_),
    .Y(_01984_));
 sky130_fd_sc_hd__mux2_1 _07957_ (.A0(_01984_),
    .A1(\LC[5] ),
    .S(_01964_),
    .X(_01985_));
 sky130_fd_sc_hd__clkbuf_1 _07958_ (.A(_01985_),
    .X(_00131_));
 sky130_fd_sc_hd__inv_2 _07959_ (.A(_01964_),
    .Y(_01986_));
 sky130_fd_sc_hd__mux2_1 _07960_ (.A0(_06280_),
    .A1(\im_reg[6] ),
    .S(_01960_),
    .X(_01987_));
 sky130_fd_sc_hd__o21ai_1 _07961_ (.A1(_01962_),
    .A2(\im_reg[6] ),
    .B1(_06279_),
    .Y(_01988_));
 sky130_fd_sc_hd__nand2_1 _07962_ (.A(_01986_),
    .B(_01988_),
    .Y(_01989_));
 sky130_fd_sc_hd__a22o_1 _07963_ (.A1(_01986_),
    .A2(_01987_),
    .B1(_01989_),
    .B2(\LC[6] ),
    .X(_00132_));
 sky130_fd_sc_hd__inv_2 _07964_ (.A(\im_reg[7] ),
    .Y(_01990_));
 sky130_fd_sc_hd__a21o_1 _07965_ (.A1(_01960_),
    .A2(_01990_),
    .B1(_06280_),
    .X(_01991_));
 sky130_fd_sc_hd__nand2_1 _07966_ (.A(_01986_),
    .B(_01991_),
    .Y(_01992_));
 sky130_fd_sc_hd__o21a_1 _07967_ (.A1(_01960_),
    .A2(_06281_),
    .B1(_01986_),
    .X(_01993_));
 sky130_fd_sc_hd__nand2_1 _07968_ (.A(_01990_),
    .B(_01960_),
    .Y(_01994_));
 sky130_fd_sc_hd__a22o_1 _07969_ (.A1(\LC[7] ),
    .A2(_01992_),
    .B1(_01993_),
    .B2(_01994_),
    .X(_00133_));
 sky130_fd_sc_hd__nor2_1 _07970_ (.A(\im_reg[8] ),
    .B(_01962_),
    .Y(_01995_));
 sky130_fd_sc_hd__a21o_1 _07971_ (.A1(_01962_),
    .A2(_06283_),
    .B1(_01964_),
    .X(_01996_));
 sky130_fd_sc_hd__o22ai_1 _07972_ (.A1(_01995_),
    .A2(_01996_),
    .B1(_06282_),
    .B2(_01993_),
    .Y(_00134_));
 sky130_fd_sc_hd__nor2_1 _07973_ (.A(\LC[9] ),
    .B(_06283_),
    .Y(_01997_));
 sky130_fd_sc_hd__mux2_1 _07974_ (.A0(_01997_),
    .A1(\im_reg[9] ),
    .S(_01960_),
    .X(_01998_));
 sky130_fd_sc_hd__a22o_1 _07975_ (.A1(_01986_),
    .A2(_01998_),
    .B1(_01996_),
    .B2(\LC[9] ),
    .X(_00135_));
 sky130_fd_sc_hd__nand2_2 _07976_ (.A(_01242_),
    .B(_01247_),
    .Y(_01999_));
 sky130_fd_sc_hd__nor2_4 _07977_ (.A(_01940_),
    .B(_01999_),
    .Y(_02000_));
 sky130_fd_sc_hd__buf_4 _07978_ (.A(_02000_),
    .X(_02001_));
 sky130_fd_sc_hd__mux2_1 _07979_ (.A0(\Oset[0][0] ),
    .A1(_01218_),
    .S(_02001_),
    .X(_02002_));
 sky130_fd_sc_hd__clkbuf_1 _07980_ (.A(_02002_),
    .X(_00136_));
 sky130_fd_sc_hd__mux2_1 _07981_ (.A0(\Oset[0][1] ),
    .A1(_01278_),
    .S(_02001_),
    .X(_02003_));
 sky130_fd_sc_hd__clkbuf_1 _07982_ (.A(_02003_),
    .X(_00137_));
 sky130_fd_sc_hd__mux2_1 _07983_ (.A0(\Oset[0][2] ),
    .A1(_01295_),
    .S(_02001_),
    .X(_02004_));
 sky130_fd_sc_hd__clkbuf_1 _07984_ (.A(_02004_),
    .X(_00138_));
 sky130_fd_sc_hd__mux2_1 _07985_ (.A0(\Oset[0][3] ),
    .A1(_01314_),
    .S(_02001_),
    .X(_02005_));
 sky130_fd_sc_hd__clkbuf_1 _07986_ (.A(_02005_),
    .X(_00139_));
 sky130_fd_sc_hd__mux2_1 _07987_ (.A0(\Oset[0][4] ),
    .A1(_01332_),
    .S(_02001_),
    .X(_02006_));
 sky130_fd_sc_hd__clkbuf_1 _07988_ (.A(_02006_),
    .X(_00140_));
 sky130_fd_sc_hd__mux2_1 _07989_ (.A0(\Oset[0][5] ),
    .A1(_01349_),
    .S(_02001_),
    .X(_02007_));
 sky130_fd_sc_hd__clkbuf_1 _07990_ (.A(_02007_),
    .X(_00141_));
 sky130_fd_sc_hd__mux2_1 _07991_ (.A0(\Oset[0][6] ),
    .A1(_01368_),
    .S(_02001_),
    .X(_02008_));
 sky130_fd_sc_hd__clkbuf_1 _07992_ (.A(_02008_),
    .X(_00142_));
 sky130_fd_sc_hd__mux2_1 _07993_ (.A0(\Oset[0][7] ),
    .A1(_01385_),
    .S(_02001_),
    .X(_02009_));
 sky130_fd_sc_hd__clkbuf_1 _07994_ (.A(_02009_),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _07995_ (.A0(\Oset[0][8] ),
    .A1(_01403_),
    .S(_02001_),
    .X(_02010_));
 sky130_fd_sc_hd__clkbuf_1 _07996_ (.A(_02010_),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _07997_ (.A0(\Oset[0][9] ),
    .A1(_01420_),
    .S(_02001_),
    .X(_02011_));
 sky130_fd_sc_hd__clkbuf_1 _07998_ (.A(_02011_),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _07999_ (.A0(\Oset[0][10] ),
    .A1(_01437_),
    .S(_02000_),
    .X(_02012_));
 sky130_fd_sc_hd__clkbuf_1 _08000_ (.A(_02012_),
    .X(_00146_));
 sky130_fd_sc_hd__mux2_1 _08001_ (.A0(\Oset[0][11] ),
    .A1(_01455_),
    .S(_02000_),
    .X(_02013_));
 sky130_fd_sc_hd__clkbuf_1 _08002_ (.A(_02013_),
    .X(_00147_));
 sky130_fd_sc_hd__mux2_1 _08003_ (.A0(\Oset[0][12] ),
    .A1(_01473_),
    .S(_02000_),
    .X(_02014_));
 sky130_fd_sc_hd__clkbuf_1 _08004_ (.A(_02014_),
    .X(_00148_));
 sky130_fd_sc_hd__mux2_1 _08005_ (.A0(\Oset[0][13] ),
    .A1(_01490_),
    .S(_02000_),
    .X(_02015_));
 sky130_fd_sc_hd__clkbuf_1 _08006_ (.A(_02015_),
    .X(_00149_));
 sky130_fd_sc_hd__mux2_1 _08007_ (.A0(\Oset[0][14] ),
    .A1(_01508_),
    .S(_02000_),
    .X(_02016_));
 sky130_fd_sc_hd__clkbuf_1 _08008_ (.A(_02016_),
    .X(_00150_));
 sky130_fd_sc_hd__mux2_1 _08009_ (.A0(\Oset[0][15] ),
    .A1(_01525_),
    .S(_02000_),
    .X(_02017_));
 sky130_fd_sc_hd__clkbuf_1 _08010_ (.A(_02017_),
    .X(_00151_));
 sky130_fd_sc_hd__nor2_4 _08011_ (.A(_01225_),
    .B(_01999_),
    .Y(_02018_));
 sky130_fd_sc_hd__buf_4 _08012_ (.A(_02018_),
    .X(_02019_));
 sky130_fd_sc_hd__mux2_1 _08013_ (.A0(\Oset[1][0] ),
    .A1(_01218_),
    .S(_02019_),
    .X(_02020_));
 sky130_fd_sc_hd__clkbuf_1 _08014_ (.A(_02020_),
    .X(_00152_));
 sky130_fd_sc_hd__mux2_1 _08015_ (.A0(\Oset[1][1] ),
    .A1(_01278_),
    .S(_02019_),
    .X(_02021_));
 sky130_fd_sc_hd__clkbuf_1 _08016_ (.A(_02021_),
    .X(_00153_));
 sky130_fd_sc_hd__mux2_1 _08017_ (.A0(\Oset[1][2] ),
    .A1(_01295_),
    .S(_02019_),
    .X(_02022_));
 sky130_fd_sc_hd__clkbuf_1 _08018_ (.A(_02022_),
    .X(_00154_));
 sky130_fd_sc_hd__mux2_1 _08019_ (.A0(\Oset[1][3] ),
    .A1(_01314_),
    .S(_02019_),
    .X(_02023_));
 sky130_fd_sc_hd__clkbuf_1 _08020_ (.A(_02023_),
    .X(_00155_));
 sky130_fd_sc_hd__mux2_1 _08021_ (.A0(\Oset[1][4] ),
    .A1(_01332_),
    .S(_02019_),
    .X(_02024_));
 sky130_fd_sc_hd__clkbuf_1 _08022_ (.A(_02024_),
    .X(_00156_));
 sky130_fd_sc_hd__mux2_1 _08023_ (.A0(\Oset[1][5] ),
    .A1(_01349_),
    .S(_02019_),
    .X(_02025_));
 sky130_fd_sc_hd__clkbuf_1 _08024_ (.A(_02025_),
    .X(_00157_));
 sky130_fd_sc_hd__mux2_1 _08025_ (.A0(\Oset[1][6] ),
    .A1(_01368_),
    .S(_02019_),
    .X(_02026_));
 sky130_fd_sc_hd__clkbuf_1 _08026_ (.A(_02026_),
    .X(_00158_));
 sky130_fd_sc_hd__mux2_1 _08027_ (.A0(\Oset[1][7] ),
    .A1(_01385_),
    .S(_02019_),
    .X(_02027_));
 sky130_fd_sc_hd__clkbuf_1 _08028_ (.A(_02027_),
    .X(_00159_));
 sky130_fd_sc_hd__mux2_1 _08029_ (.A0(\Oset[1][8] ),
    .A1(_01403_),
    .S(_02019_),
    .X(_02028_));
 sky130_fd_sc_hd__clkbuf_1 _08030_ (.A(_02028_),
    .X(_00160_));
 sky130_fd_sc_hd__mux2_1 _08031_ (.A0(\Oset[1][9] ),
    .A1(_01420_),
    .S(_02019_),
    .X(_02029_));
 sky130_fd_sc_hd__clkbuf_1 _08032_ (.A(_02029_),
    .X(_00161_));
 sky130_fd_sc_hd__mux2_1 _08033_ (.A0(\Oset[1][10] ),
    .A1(_01437_),
    .S(_02018_),
    .X(_02030_));
 sky130_fd_sc_hd__clkbuf_1 _08034_ (.A(_02030_),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _08035_ (.A0(\Oset[1][11] ),
    .A1(_01455_),
    .S(_02018_),
    .X(_02031_));
 sky130_fd_sc_hd__clkbuf_1 _08036_ (.A(_02031_),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _08037_ (.A0(\Oset[1][12] ),
    .A1(_01473_),
    .S(_02018_),
    .X(_02032_));
 sky130_fd_sc_hd__clkbuf_1 _08038_ (.A(_02032_),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _08039_ (.A0(\Oset[1][13] ),
    .A1(_01490_),
    .S(_02018_),
    .X(_02033_));
 sky130_fd_sc_hd__clkbuf_1 _08040_ (.A(_02033_),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _08041_ (.A0(\Oset[1][14] ),
    .A1(_01508_),
    .S(_02018_),
    .X(_02034_));
 sky130_fd_sc_hd__clkbuf_1 _08042_ (.A(_02034_),
    .X(_00166_));
 sky130_fd_sc_hd__mux2_1 _08043_ (.A0(\Oset[1][15] ),
    .A1(_01525_),
    .S(_02018_),
    .X(_02035_));
 sky130_fd_sc_hd__clkbuf_1 _08044_ (.A(_02035_),
    .X(_00167_));
 sky130_fd_sc_hd__or2_1 _08045_ (.A(_01627_),
    .B(_01623_),
    .X(_02036_));
 sky130_fd_sc_hd__clkbuf_4 _08046_ (.A(_02036_),
    .X(_02037_));
 sky130_fd_sc_hd__clkbuf_8 _08047_ (.A(_02037_),
    .X(_02038_));
 sky130_fd_sc_hd__mux2_1 _08048_ (.A0(_01615_),
    .A1(\H[2][0] ),
    .S(_02038_),
    .X(_02039_));
 sky130_fd_sc_hd__clkbuf_1 _08049_ (.A(_02039_),
    .X(_00168_));
 sky130_fd_sc_hd__mux2_1 _08050_ (.A0(_01650_),
    .A1(\H[2][1] ),
    .S(_02038_),
    .X(_02040_));
 sky130_fd_sc_hd__clkbuf_1 _08051_ (.A(_02040_),
    .X(_00169_));
 sky130_fd_sc_hd__mux2_1 _08052_ (.A0(_01676_),
    .A1(\H[2][2] ),
    .S(_02038_),
    .X(_02041_));
 sky130_fd_sc_hd__clkbuf_1 _08053_ (.A(_02041_),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _08054_ (.A0(_01700_),
    .A1(\H[2][3] ),
    .S(_02038_),
    .X(_02042_));
 sky130_fd_sc_hd__clkbuf_1 _08055_ (.A(_02042_),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_1 _08056_ (.A0(_01720_),
    .A1(\H[2][4] ),
    .S(_02038_),
    .X(_02043_));
 sky130_fd_sc_hd__clkbuf_1 _08057_ (.A(_02043_),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _08058_ (.A0(_01740_),
    .A1(\H[2][5] ),
    .S(_02038_),
    .X(_02044_));
 sky130_fd_sc_hd__clkbuf_1 _08059_ (.A(_02044_),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _08060_ (.A0(_01761_),
    .A1(\H[2][6] ),
    .S(_02038_),
    .X(_02045_));
 sky130_fd_sc_hd__clkbuf_1 _08061_ (.A(_02045_),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_1 _08062_ (.A0(_01781_),
    .A1(\H[2][7] ),
    .S(_02038_),
    .X(_02046_));
 sky130_fd_sc_hd__clkbuf_1 _08063_ (.A(_02046_),
    .X(_00175_));
 sky130_fd_sc_hd__mux2_1 _08064_ (.A0(_01801_),
    .A1(\H[2][8] ),
    .S(_02038_),
    .X(_02047_));
 sky130_fd_sc_hd__clkbuf_1 _08065_ (.A(_02047_),
    .X(_00176_));
 sky130_fd_sc_hd__mux2_1 _08066_ (.A0(_01819_),
    .A1(\H[2][9] ),
    .S(_02038_),
    .X(_02048_));
 sky130_fd_sc_hd__clkbuf_1 _08067_ (.A(_02048_),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _08068_ (.A0(_01839_),
    .A1(\H[2][10] ),
    .S(_02037_),
    .X(_02049_));
 sky130_fd_sc_hd__clkbuf_1 _08069_ (.A(_02049_),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _08070_ (.A0(_01859_),
    .A1(\H[2][11] ),
    .S(_02037_),
    .X(_02050_));
 sky130_fd_sc_hd__clkbuf_1 _08071_ (.A(_02050_),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _08072_ (.A0(_01879_),
    .A1(\H[2][12] ),
    .S(_02037_),
    .X(_02051_));
 sky130_fd_sc_hd__clkbuf_1 _08073_ (.A(_02051_),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _08074_ (.A0(_01898_),
    .A1(\H[2][13] ),
    .S(_02037_),
    .X(_02052_));
 sky130_fd_sc_hd__clkbuf_1 _08075_ (.A(_02052_),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _08076_ (.A0(_01918_),
    .A1(\H[2][14] ),
    .S(_02037_),
    .X(_02053_));
 sky130_fd_sc_hd__clkbuf_1 _08077_ (.A(_02053_),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _08078_ (.A0(_01938_),
    .A1(\H[2][15] ),
    .S(_02037_),
    .X(_02054_));
 sky130_fd_sc_hd__clkbuf_1 _08079_ (.A(_02054_),
    .X(_00183_));
 sky130_fd_sc_hd__nand2_1 _08080_ (.A(_01619_),
    .B(_01622_),
    .Y(_02055_));
 sky130_fd_sc_hd__nand2b_4 _08081_ (.A_N(_02055_),
    .B(_01627_),
    .Y(_02056_));
 sky130_fd_sc_hd__buf_4 _08082_ (.A(_02056_),
    .X(_02057_));
 sky130_fd_sc_hd__mux2_1 _08083_ (.A0(_01615_),
    .A1(\H[1][0] ),
    .S(_02057_),
    .X(_02058_));
 sky130_fd_sc_hd__clkbuf_1 _08084_ (.A(_02058_),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _08085_ (.A0(_01650_),
    .A1(\H[1][1] ),
    .S(_02057_),
    .X(_02059_));
 sky130_fd_sc_hd__clkbuf_1 _08086_ (.A(_02059_),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _08087_ (.A0(_01676_),
    .A1(\H[1][2] ),
    .S(_02057_),
    .X(_02060_));
 sky130_fd_sc_hd__clkbuf_1 _08088_ (.A(_02060_),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _08089_ (.A0(_01700_),
    .A1(\H[1][3] ),
    .S(_02057_),
    .X(_02061_));
 sky130_fd_sc_hd__clkbuf_1 _08090_ (.A(_02061_),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _08091_ (.A0(_01720_),
    .A1(\H[1][4] ),
    .S(_02057_),
    .X(_02062_));
 sky130_fd_sc_hd__clkbuf_1 _08092_ (.A(_02062_),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _08093_ (.A0(_01740_),
    .A1(\H[1][5] ),
    .S(_02057_),
    .X(_02063_));
 sky130_fd_sc_hd__clkbuf_1 _08094_ (.A(_02063_),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _08095_ (.A0(_01761_),
    .A1(\H[1][6] ),
    .S(_02057_),
    .X(_02064_));
 sky130_fd_sc_hd__clkbuf_1 _08096_ (.A(_02064_),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _08097_ (.A0(_01781_),
    .A1(\H[1][7] ),
    .S(_02057_),
    .X(_02065_));
 sky130_fd_sc_hd__clkbuf_1 _08098_ (.A(_02065_),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _08099_ (.A0(_01801_),
    .A1(\H[1][8] ),
    .S(_02057_),
    .X(_02066_));
 sky130_fd_sc_hd__clkbuf_1 _08100_ (.A(_02066_),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _08101_ (.A0(_01819_),
    .A1(\H[1][9] ),
    .S(_02057_),
    .X(_02067_));
 sky130_fd_sc_hd__clkbuf_1 _08102_ (.A(_02067_),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _08103_ (.A0(_01839_),
    .A1(\H[1][10] ),
    .S(_02056_),
    .X(_02068_));
 sky130_fd_sc_hd__clkbuf_1 _08104_ (.A(_02068_),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _08105_ (.A0(_01859_),
    .A1(\H[1][11] ),
    .S(_02056_),
    .X(_02069_));
 sky130_fd_sc_hd__clkbuf_1 _08106_ (.A(_02069_),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_1 _08107_ (.A0(_01879_),
    .A1(\H[1][12] ),
    .S(_02056_),
    .X(_02070_));
 sky130_fd_sc_hd__clkbuf_1 _08108_ (.A(_02070_),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _08109_ (.A0(_01898_),
    .A1(\H[1][13] ),
    .S(_02056_),
    .X(_02071_));
 sky130_fd_sc_hd__clkbuf_1 _08110_ (.A(_02071_),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _08111_ (.A0(_01918_),
    .A1(\H[1][14] ),
    .S(_02056_),
    .X(_02072_));
 sky130_fd_sc_hd__clkbuf_1 _08112_ (.A(_02072_),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _08113_ (.A0(_01938_),
    .A1(\H[1][15] ),
    .S(_02056_),
    .X(_02073_));
 sky130_fd_sc_hd__clkbuf_1 _08114_ (.A(_02073_),
    .X(_00199_));
 sky130_fd_sc_hd__nor2_4 _08115_ (.A(_01627_),
    .B(_02055_),
    .Y(_02074_));
 sky130_fd_sc_hd__clkbuf_8 _08116_ (.A(_02074_),
    .X(_02075_));
 sky130_fd_sc_hd__mux2_1 _08117_ (.A0(\H[0][0] ),
    .A1(_01615_),
    .S(_02075_),
    .X(_02076_));
 sky130_fd_sc_hd__clkbuf_1 _08118_ (.A(_02076_),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _08119_ (.A0(\H[0][1] ),
    .A1(_01650_),
    .S(_02075_),
    .X(_02077_));
 sky130_fd_sc_hd__clkbuf_1 _08120_ (.A(_02077_),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _08121_ (.A0(\H[0][2] ),
    .A1(_01676_),
    .S(_02075_),
    .X(_02078_));
 sky130_fd_sc_hd__clkbuf_1 _08122_ (.A(_02078_),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _08123_ (.A0(\H[0][3] ),
    .A1(_01700_),
    .S(_02075_),
    .X(_02079_));
 sky130_fd_sc_hd__clkbuf_1 _08124_ (.A(_02079_),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _08125_ (.A0(\H[0][4] ),
    .A1(_01720_),
    .S(_02075_),
    .X(_02080_));
 sky130_fd_sc_hd__clkbuf_1 _08126_ (.A(_02080_),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _08127_ (.A0(\H[0][5] ),
    .A1(_01740_),
    .S(_02075_),
    .X(_02081_));
 sky130_fd_sc_hd__clkbuf_1 _08128_ (.A(_02081_),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _08129_ (.A0(\H[0][6] ),
    .A1(_01761_),
    .S(_02075_),
    .X(_02082_));
 sky130_fd_sc_hd__clkbuf_1 _08130_ (.A(_02082_),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_1 _08131_ (.A0(\H[0][7] ),
    .A1(_01781_),
    .S(_02075_),
    .X(_02083_));
 sky130_fd_sc_hd__clkbuf_1 _08132_ (.A(_02083_),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _08133_ (.A0(\H[0][8] ),
    .A1(_01801_),
    .S(_02075_),
    .X(_02084_));
 sky130_fd_sc_hd__clkbuf_1 _08134_ (.A(_02084_),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _08135_ (.A0(\H[0][9] ),
    .A1(_01819_),
    .S(_02075_),
    .X(_02085_));
 sky130_fd_sc_hd__clkbuf_1 _08136_ (.A(_02085_),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _08137_ (.A0(\H[0][10] ),
    .A1(_01839_),
    .S(_02074_),
    .X(_02086_));
 sky130_fd_sc_hd__clkbuf_1 _08138_ (.A(_02086_),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _08139_ (.A0(\H[0][11] ),
    .A1(_01859_),
    .S(_02074_),
    .X(_02087_));
 sky130_fd_sc_hd__clkbuf_1 _08140_ (.A(_02087_),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _08141_ (.A0(\H[0][12] ),
    .A1(_01879_),
    .S(_02074_),
    .X(_02088_));
 sky130_fd_sc_hd__clkbuf_1 _08142_ (.A(_02088_),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _08143_ (.A0(\H[0][13] ),
    .A1(_01898_),
    .S(_02074_),
    .X(_02089_));
 sky130_fd_sc_hd__clkbuf_1 _08144_ (.A(_02089_),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _08145_ (.A0(\H[0][14] ),
    .A1(_01918_),
    .S(_02074_),
    .X(_02090_));
 sky130_fd_sc_hd__clkbuf_1 _08146_ (.A(_02090_),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _08147_ (.A0(\H[0][15] ),
    .A1(_01938_),
    .S(_02074_),
    .X(_02091_));
 sky130_fd_sc_hd__clkbuf_1 _08148_ (.A(_02091_),
    .X(_00215_));
 sky130_fd_sc_hd__clkbuf_4 _08149_ (.A(\Add.sub ),
    .X(_02092_));
 sky130_fd_sc_hd__nor2_1 _08150_ (.A(_02092_),
    .B(CMD_addition),
    .Y(_02093_));
 sky130_fd_sc_hd__o211a_1 _08151_ (.A1(CMD_store),
    .A2(CMD_load),
    .B1(_00597_),
    .C1(_02093_),
    .X(_02094_));
 sky130_fd_sc_hd__and3_2 _08152_ (.A(_02094_),
    .B(_00578_),
    .C(_00546_),
    .X(_02095_));
 sky130_fd_sc_hd__buf_4 _08153_ (.A(_00556_),
    .X(_02096_));
 sky130_fd_sc_hd__and3_1 _08154_ (.A(_00547_),
    .B(_02096_),
    .C(\current_state[6] ),
    .X(_02097_));
 sky130_fd_sc_hd__inv_2 _08155_ (.A(_02097_),
    .Y(_02098_));
 sky130_fd_sc_hd__nor2_4 _08156_ (.A(_00557_),
    .B(_02098_),
    .Y(_02099_));
 sky130_fd_sc_hd__nand2_4 _08157_ (.A(_02095_),
    .B(_02099_),
    .Y(_02100_));
 sky130_fd_sc_hd__buf_4 _08158_ (.A(_01148_),
    .X(_02101_));
 sky130_fd_sc_hd__buf_2 _08159_ (.A(_02095_),
    .X(_02102_));
 sky130_fd_sc_hd__buf_2 _08160_ (.A(_02099_),
    .X(_02103_));
 sky130_fd_sc_hd__a21o_1 _08161_ (.A1(_02102_),
    .A2(_02103_),
    .B1(net38),
    .X(_02104_));
 sky130_fd_sc_hd__o211a_1 _08162_ (.A1(\R3[0] ),
    .A2(_02100_),
    .B1(_02101_),
    .C1(_02104_),
    .X(_00216_));
 sky130_fd_sc_hd__buf_4 _08163_ (.A(_01148_),
    .X(_02105_));
 sky130_fd_sc_hd__a21o_1 _08164_ (.A1(_02102_),
    .A2(_02103_),
    .B1(net39),
    .X(_02106_));
 sky130_fd_sc_hd__o211a_1 _08165_ (.A1(\R3[1] ),
    .A2(_02100_),
    .B1(_02105_),
    .C1(_02106_),
    .X(_00217_));
 sky130_fd_sc_hd__a21o_1 _08166_ (.A1(_02102_),
    .A2(_02103_),
    .B1(net40),
    .X(_02107_));
 sky130_fd_sc_hd__o211a_1 _08167_ (.A1(\R2[0] ),
    .A2(_02100_),
    .B1(_02105_),
    .C1(_02107_),
    .X(_00218_));
 sky130_fd_sc_hd__a21o_1 _08168_ (.A1(_02102_),
    .A2(_02103_),
    .B1(net41),
    .X(_02108_));
 sky130_fd_sc_hd__o211a_1 _08169_ (.A1(\R2[1] ),
    .A2(_02100_),
    .B1(_02105_),
    .C1(_02108_),
    .X(_00219_));
 sky130_fd_sc_hd__a21o_1 _08170_ (.A1(_02102_),
    .A2(_02103_),
    .B1(net42),
    .X(_02109_));
 sky130_fd_sc_hd__o211a_1 _08171_ (.A1(_00498_),
    .A2(_02100_),
    .B1(_02105_),
    .C1(_02109_),
    .X(_00220_));
 sky130_fd_sc_hd__a21o_1 _08172_ (.A1(_02102_),
    .A2(_02103_),
    .B1(net43),
    .X(_02110_));
 sky130_fd_sc_hd__o211a_1 _08173_ (.A1(\R1[1] ),
    .A2(_02100_),
    .B1(_02105_),
    .C1(_02110_),
    .X(_00221_));
 sky130_fd_sc_hd__a21o_1 _08174_ (.A1(_02102_),
    .A2(_02103_),
    .B1(net44),
    .X(_02111_));
 sky130_fd_sc_hd__o211a_1 _08175_ (.A1(\im_reg[6] ),
    .A2(_02100_),
    .B1(_02105_),
    .C1(_02111_),
    .X(_00222_));
 sky130_fd_sc_hd__a21o_1 _08176_ (.A1(_02102_),
    .A2(_02103_),
    .B1(net45),
    .X(_02112_));
 sky130_fd_sc_hd__o211a_1 _08177_ (.A1(\im_reg[7] ),
    .A2(_02100_),
    .B1(_02105_),
    .C1(_02112_),
    .X(_00223_));
 sky130_fd_sc_hd__a21o_1 _08178_ (.A1(_02102_),
    .A2(_02103_),
    .B1(net46),
    .X(_02113_));
 sky130_fd_sc_hd__o211a_1 _08179_ (.A1(\im_reg[8] ),
    .A2(_02100_),
    .B1(_02105_),
    .C1(_02113_),
    .X(_00224_));
 sky130_fd_sc_hd__a21o_1 _08180_ (.A1(_02095_),
    .A2(_02099_),
    .B1(net47),
    .X(_02114_));
 sky130_fd_sc_hd__o211a_1 _08181_ (.A1(\im_reg[9] ),
    .A2(_02100_),
    .B1(_02105_),
    .C1(_02114_),
    .X(_00225_));
 sky130_fd_sc_hd__buf_4 _08182_ (.A(_00635_),
    .X(_02115_));
 sky130_fd_sc_hd__buf_4 _08183_ (.A(_02115_),
    .X(_02116_));
 sky130_fd_sc_hd__a21oi_1 _08184_ (.A1(_02102_),
    .A2(_02103_),
    .B1(net36),
    .Y(_02117_));
 sky130_fd_sc_hd__nor2_1 _08185_ (.A(_02116_),
    .B(_02117_),
    .Y(_00226_));
 sky130_fd_sc_hd__buf_4 _08186_ (.A(\shift.left ),
    .X(_02118_));
 sky130_fd_sc_hd__nor2_1 _08187_ (.A(_02118_),
    .B(CMD_addition),
    .Y(_02119_));
 sky130_fd_sc_hd__nor2_1 _08188_ (.A(CMD_not),
    .B(CMD_logic_shift_right),
    .Y(_02120_));
 sky130_fd_sc_hd__nand2_1 _08189_ (.A(_02119_),
    .B(_02120_),
    .Y(_02121_));
 sky130_fd_sc_hd__nand3_1 _08190_ (.A(_00597_),
    .B(CMD_store),
    .C(_00697_),
    .Y(_02122_));
 sky130_fd_sc_hd__nor2_1 _08191_ (.A(_02121_),
    .B(_02122_),
    .Y(_02123_));
 sky130_fd_sc_hd__and3_1 _08192_ (.A(_02123_),
    .B(_00832_),
    .C(_02099_),
    .X(_02124_));
 sky130_fd_sc_hd__buf_4 _08193_ (.A(_01148_),
    .X(_02125_));
 sky130_fd_sc_hd__o21a_1 _08194_ (.A1(net37),
    .A2(_02124_),
    .B1(_02125_),
    .X(_00227_));
 sky130_fd_sc_hd__buf_8 _08195_ (.A(_00591_),
    .X(_02126_));
 sky130_fd_sc_hd__buf_6 _08196_ (.A(_00002_),
    .X(_02127_));
 sky130_fd_sc_hd__inv_6 _08197_ (.A(_02127_),
    .Y(_02128_));
 sky130_fd_sc_hd__buf_6 _08198_ (.A(_02128_),
    .X(_02129_));
 sky130_fd_sc_hd__nand2_1 _08199_ (.A(_02129_),
    .B(\Qset[2][0] ),
    .Y(_02130_));
 sky130_fd_sc_hd__buf_4 _08200_ (.A(_02127_),
    .X(_02131_));
 sky130_fd_sc_hd__nand2_1 _08201_ (.A(\Qset[3][0] ),
    .B(_02131_),
    .Y(_02132_));
 sky130_fd_sc_hd__nand3_1 _08202_ (.A(_02130_),
    .B(_00003_),
    .C(_02132_),
    .Y(_02133_));
 sky130_fd_sc_hd__nand2_1 _08203_ (.A(_02129_),
    .B(\Qset[0][0] ),
    .Y(_02134_));
 sky130_fd_sc_hd__inv_2 _08204_ (.A(_00003_),
    .Y(_02135_));
 sky130_fd_sc_hd__nand2_1 _08205_ (.A(\Qset[1][0] ),
    .B(_02131_),
    .Y(_02136_));
 sky130_fd_sc_hd__nand3_1 _08206_ (.A(_02134_),
    .B(_02135_),
    .C(_02136_),
    .Y(_02137_));
 sky130_fd_sc_hd__nand2_1 _08207_ (.A(_02133_),
    .B(_02137_),
    .Y(_02138_));
 sky130_fd_sc_hd__buf_8 _08208_ (.A(_01162_),
    .X(_02139_));
 sky130_fd_sc_hd__buf_8 _08209_ (.A(_02139_),
    .X(_02140_));
 sky130_fd_sc_hd__buf_6 _08210_ (.A(_02127_),
    .X(_02141_));
 sky130_fd_sc_hd__inv_2 _08211_ (.A(\Oset[2][0] ),
    .Y(_02142_));
 sky130_fd_sc_hd__clkbuf_4 _08212_ (.A(_00003_),
    .X(_02143_));
 sky130_fd_sc_hd__nand2_1 _08213_ (.A(_02141_),
    .B(\Oset[3][0] ),
    .Y(_02144_));
 sky130_fd_sc_hd__o211ai_1 _08214_ (.A1(_02141_),
    .A2(_02142_),
    .B1(_02143_),
    .C1(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__inv_2 _08215_ (.A(\Oset[0][0] ),
    .Y(_02146_));
 sky130_fd_sc_hd__buf_4 _08216_ (.A(_02135_),
    .X(_02147_));
 sky130_fd_sc_hd__nand2_1 _08217_ (.A(_02141_),
    .B(\Oset[1][0] ),
    .Y(_02148_));
 sky130_fd_sc_hd__o211ai_1 _08218_ (.A1(_02131_),
    .A2(_02146_),
    .B1(_02147_),
    .C1(_02148_),
    .Y(_02149_));
 sky130_fd_sc_hd__nand2_1 _08219_ (.A(_02145_),
    .B(_02149_),
    .Y(_02150_));
 sky130_fd_sc_hd__buf_2 _08220_ (.A(_02128_),
    .X(_02151_));
 sky130_fd_sc_hd__inv_2 _08221_ (.A(\H[2][0] ),
    .Y(_02152_));
 sky130_fd_sc_hd__nor2_1 _08222_ (.A(\H[3][0] ),
    .B(_02151_),
    .Y(_02153_));
 sky130_fd_sc_hd__a211o_1 _08223_ (.A1(_02151_),
    .A2(_02152_),
    .B1(_02147_),
    .C1(_02153_),
    .X(_02154_));
 sky130_fd_sc_hd__inv_2 _08224_ (.A(\H[0][0] ),
    .Y(_02155_));
 sky130_fd_sc_hd__nor2_1 _08225_ (.A(\H[1][0] ),
    .B(_02151_),
    .Y(_02156_));
 sky130_fd_sc_hd__a211o_1 _08226_ (.A1(_02151_),
    .A2(_02155_),
    .B1(_02143_),
    .C1(_02156_),
    .X(_02157_));
 sky130_fd_sc_hd__a21o_2 _08227_ (.A1(_02154_),
    .A2(_02157_),
    .B1(_01551_),
    .X(_02158_));
 sky130_fd_sc_hd__o221ai_4 _08228_ (.A1(_02126_),
    .A2(_02138_),
    .B1(_02140_),
    .B2(_02150_),
    .C1(_02158_),
    .Y(_02159_));
 sky130_fd_sc_hd__buf_4 _08229_ (.A(_02092_),
    .X(_02160_));
 sky130_fd_sc_hd__clkbuf_4 _08230_ (.A(\shift.Q ),
    .X(_02161_));
 sky130_fd_sc_hd__clkbuf_4 _08231_ (.A(_02161_),
    .X(_02162_));
 sky130_fd_sc_hd__clkbuf_4 _08232_ (.A(_02162_),
    .X(_02163_));
 sky130_fd_sc_hd__nor2_1 _08233_ (.A(_02163_),
    .B(_00591_),
    .Y(_02164_));
 sky130_fd_sc_hd__nor2_1 _08234_ (.A(_02160_),
    .B(_02164_),
    .Y(_02165_));
 sky130_fd_sc_hd__nand2_1 _08235_ (.A(_02165_),
    .B(_02123_),
    .Y(_02166_));
 sky130_fd_sc_hd__inv_2 _08236_ (.A(_02099_),
    .Y(_02167_));
 sky130_fd_sc_hd__or3_2 _08237_ (.A(_00635_),
    .B(_02166_),
    .C(_02167_),
    .X(_02168_));
 sky130_fd_sc_hd__clkbuf_4 _08238_ (.A(_02168_),
    .X(_02169_));
 sky130_fd_sc_hd__clkbuf_4 _08239_ (.A(_02169_),
    .X(_02170_));
 sky130_fd_sc_hd__mux2_1 _08240_ (.A0(_02159_),
    .A1(net48),
    .S(_02170_),
    .X(_02171_));
 sky130_fd_sc_hd__clkbuf_1 _08241_ (.A(_02171_),
    .X(_00228_));
 sky130_fd_sc_hd__nand2_1 _08242_ (.A(_02128_),
    .B(\Qset[2][1] ),
    .Y(_02172_));
 sky130_fd_sc_hd__nand2_1 _08243_ (.A(_02127_),
    .B(\Qset[3][1] ),
    .Y(_02173_));
 sky130_fd_sc_hd__nand3_1 _08244_ (.A(_02172_),
    .B(_00003_),
    .C(_02173_),
    .Y(_02174_));
 sky130_fd_sc_hd__nand2_1 _08245_ (.A(_02128_),
    .B(\Qset[0][1] ),
    .Y(_02175_));
 sky130_fd_sc_hd__nand2_1 _08246_ (.A(_02127_),
    .B(\Qset[1][1] ),
    .Y(_02176_));
 sky130_fd_sc_hd__nand3_1 _08247_ (.A(_02175_),
    .B(_02135_),
    .C(_02176_),
    .Y(_02177_));
 sky130_fd_sc_hd__nand2_2 _08248_ (.A(_02174_),
    .B(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__inv_2 _08249_ (.A(\Oset[2][1] ),
    .Y(_02179_));
 sky130_fd_sc_hd__nand2_1 _08250_ (.A(_02131_),
    .B(\Oset[3][1] ),
    .Y(_02180_));
 sky130_fd_sc_hd__o211ai_1 _08251_ (.A1(_02131_),
    .A2(_02179_),
    .B1(_00003_),
    .C1(_02180_),
    .Y(_02181_));
 sky130_fd_sc_hd__inv_2 _08252_ (.A(\Oset[0][1] ),
    .Y(_02182_));
 sky130_fd_sc_hd__nand2_1 _08253_ (.A(_02127_),
    .B(\Oset[1][1] ),
    .Y(_02183_));
 sky130_fd_sc_hd__o211ai_1 _08254_ (.A1(_02127_),
    .A2(_02182_),
    .B1(_02135_),
    .C1(_02183_),
    .Y(_02184_));
 sky130_fd_sc_hd__nand2_1 _08255_ (.A(_02181_),
    .B(_02184_),
    .Y(_02185_));
 sky130_fd_sc_hd__inv_2 _08256_ (.A(\H[2][1] ),
    .Y(_02186_));
 sky130_fd_sc_hd__nor2_1 _08257_ (.A(\H[3][1] ),
    .B(_02129_),
    .Y(_02187_));
 sky130_fd_sc_hd__a211o_1 _08258_ (.A1(_02129_),
    .A2(_02186_),
    .B1(_02135_),
    .C1(_02187_),
    .X(_02188_));
 sky130_fd_sc_hd__inv_2 _08259_ (.A(\H[0][1] ),
    .Y(_02189_));
 sky130_fd_sc_hd__nor2_1 _08260_ (.A(\H[1][1] ),
    .B(_02129_),
    .Y(_02190_));
 sky130_fd_sc_hd__a211o_1 _08261_ (.A1(_02129_),
    .A2(_02189_),
    .B1(_00003_),
    .C1(_02190_),
    .X(_02191_));
 sky130_fd_sc_hd__a21o_1 _08262_ (.A1(_02188_),
    .A2(_02191_),
    .B1(_01551_),
    .X(_02192_));
 sky130_fd_sc_hd__o221ai_2 _08263_ (.A1(_02126_),
    .A2(_02178_),
    .B1(_02140_),
    .B2(_02185_),
    .C1(_02192_),
    .Y(_02193_));
 sky130_fd_sc_hd__mux2_1 _08264_ (.A0(_02193_),
    .A1(net55),
    .S(_02170_),
    .X(_02194_));
 sky130_fd_sc_hd__clkbuf_1 _08265_ (.A(_02194_),
    .X(_00229_));
 sky130_fd_sc_hd__nand2_1 _08266_ (.A(_02128_),
    .B(\Qset[2][2] ),
    .Y(_02195_));
 sky130_fd_sc_hd__nand2_1 _08267_ (.A(_02127_),
    .B(\Qset[3][2] ),
    .Y(_02196_));
 sky130_fd_sc_hd__nand3_1 _08268_ (.A(_02195_),
    .B(_00003_),
    .C(_02196_),
    .Y(_02197_));
 sky130_fd_sc_hd__nand2_1 _08269_ (.A(_02128_),
    .B(\Qset[0][2] ),
    .Y(_02198_));
 sky130_fd_sc_hd__nand2_1 _08270_ (.A(_02127_),
    .B(\Qset[1][2] ),
    .Y(_02199_));
 sky130_fd_sc_hd__nand3_1 _08271_ (.A(_02198_),
    .B(_02135_),
    .C(_02199_),
    .Y(_02200_));
 sky130_fd_sc_hd__nand2_1 _08272_ (.A(_02197_),
    .B(_02200_),
    .Y(_02201_));
 sky130_fd_sc_hd__nor2_1 _08273_ (.A(\Oset[3][2] ),
    .B(_02129_),
    .Y(_02202_));
 sky130_fd_sc_hd__o21ai_1 _08274_ (.A1(_02127_),
    .A2(\Oset[2][2] ),
    .B1(_00003_),
    .Y(_02203_));
 sky130_fd_sc_hd__nor2_1 _08275_ (.A(_02131_),
    .B(\Oset[0][2] ),
    .Y(_02204_));
 sky130_fd_sc_hd__o21ai_1 _08276_ (.A1(\Oset[1][2] ),
    .A2(_02129_),
    .B1(_02135_),
    .Y(_02205_));
 sky130_fd_sc_hd__o22a_1 _08277_ (.A1(_02202_),
    .A2(_02203_),
    .B1(_02204_),
    .B2(_02205_),
    .X(_02206_));
 sky130_fd_sc_hd__inv_2 _08278_ (.A(\H[2][2] ),
    .Y(_02207_));
 sky130_fd_sc_hd__nor2_1 _08279_ (.A(\H[3][2] ),
    .B(_02151_),
    .Y(_02208_));
 sky130_fd_sc_hd__a211o_1 _08280_ (.A1(_02151_),
    .A2(_02207_),
    .B1(_02147_),
    .C1(_02208_),
    .X(_02209_));
 sky130_fd_sc_hd__inv_2 _08281_ (.A(\H[0][2] ),
    .Y(_02210_));
 sky130_fd_sc_hd__nor2_1 _08282_ (.A(\H[1][2] ),
    .B(_02129_),
    .Y(_02211_));
 sky130_fd_sc_hd__a211o_1 _08283_ (.A1(_02151_),
    .A2(_02210_),
    .B1(_00003_),
    .C1(_02211_),
    .X(_02212_));
 sky130_fd_sc_hd__a21o_1 _08284_ (.A1(_02209_),
    .A2(_02212_),
    .B1(_01551_),
    .X(_02213_));
 sky130_fd_sc_hd__o221ai_2 _08285_ (.A1(_02126_),
    .A2(_02201_),
    .B1(_02140_),
    .B2(_02206_),
    .C1(_02213_),
    .Y(_02214_));
 sky130_fd_sc_hd__mux2_1 _08286_ (.A0(_02214_),
    .A1(net56),
    .S(_02170_),
    .X(_02215_));
 sky130_fd_sc_hd__clkbuf_1 _08287_ (.A(_02215_),
    .X(_00230_));
 sky130_fd_sc_hd__nand2_1 _08288_ (.A(_02151_),
    .B(\Qset[2][3] ),
    .Y(_02216_));
 sky130_fd_sc_hd__nand2_1 _08289_ (.A(_02131_),
    .B(\Qset[3][3] ),
    .Y(_02217_));
 sky130_fd_sc_hd__nand3_1 _08290_ (.A(_02216_),
    .B(_02143_),
    .C(_02217_),
    .Y(_02218_));
 sky130_fd_sc_hd__nand2_1 _08291_ (.A(_02151_),
    .B(\Qset[0][3] ),
    .Y(_02219_));
 sky130_fd_sc_hd__nand2_1 _08292_ (.A(_02131_),
    .B(\Qset[1][3] ),
    .Y(_02220_));
 sky130_fd_sc_hd__nand3_1 _08293_ (.A(_02219_),
    .B(_02147_),
    .C(_02220_),
    .Y(_02221_));
 sky130_fd_sc_hd__nand2_2 _08294_ (.A(_02218_),
    .B(_02221_),
    .Y(_02222_));
 sky130_fd_sc_hd__nand2_1 _08295_ (.A(_02131_),
    .B(\Oset[3][3] ),
    .Y(_02223_));
 sky130_fd_sc_hd__nand2_1 _08296_ (.A(_02223_),
    .B(_02143_),
    .Y(_02224_));
 sky130_fd_sc_hd__a21o_1 _08297_ (.A1(_02151_),
    .A2(\Oset[2][3] ),
    .B1(_02224_),
    .X(_02225_));
 sky130_fd_sc_hd__inv_2 _08298_ (.A(\Oset[0][3] ),
    .Y(_02226_));
 sky130_fd_sc_hd__nand2_1 _08299_ (.A(_02141_),
    .B(\Oset[1][3] ),
    .Y(_02227_));
 sky130_fd_sc_hd__o211ai_1 _08300_ (.A1(_02141_),
    .A2(_02226_),
    .B1(_02147_),
    .C1(_02227_),
    .Y(_02228_));
 sky130_fd_sc_hd__nand2_1 _08301_ (.A(_02225_),
    .B(_02228_),
    .Y(_02229_));
 sky130_fd_sc_hd__buf_6 _08302_ (.A(_02129_),
    .X(_02230_));
 sky130_fd_sc_hd__inv_2 _08303_ (.A(\H[2][3] ),
    .Y(_02231_));
 sky130_fd_sc_hd__nor2_1 _08304_ (.A(\H[3][3] ),
    .B(_02230_),
    .Y(_02232_));
 sky130_fd_sc_hd__a211o_1 _08305_ (.A1(_02230_),
    .A2(_02231_),
    .B1(_02147_),
    .C1(_02232_),
    .X(_02233_));
 sky130_fd_sc_hd__inv_2 _08306_ (.A(\H[0][3] ),
    .Y(_02234_));
 sky130_fd_sc_hd__nor2_1 _08307_ (.A(\H[1][3] ),
    .B(_02230_),
    .Y(_02235_));
 sky130_fd_sc_hd__a211o_1 _08308_ (.A1(_02230_),
    .A2(_02234_),
    .B1(_02143_),
    .C1(_02235_),
    .X(_02236_));
 sky130_fd_sc_hd__a21o_1 _08309_ (.A1(_02233_),
    .A2(_02236_),
    .B1(_01551_),
    .X(_02237_));
 sky130_fd_sc_hd__o221ai_4 _08310_ (.A1(_02126_),
    .A2(_02222_),
    .B1(_02140_),
    .B2(_02229_),
    .C1(_02237_),
    .Y(_02238_));
 sky130_fd_sc_hd__mux2_1 _08311_ (.A0(_02238_),
    .A1(net57),
    .S(_02170_),
    .X(_02239_));
 sky130_fd_sc_hd__clkbuf_1 _08312_ (.A(_02239_),
    .X(_00231_));
 sky130_fd_sc_hd__nand2_1 _08313_ (.A(_02230_),
    .B(\Qset[2][4] ),
    .Y(_02240_));
 sky130_fd_sc_hd__buf_6 _08314_ (.A(_02131_),
    .X(_02241_));
 sky130_fd_sc_hd__nand2_1 _08315_ (.A(_02241_),
    .B(\Qset[3][4] ),
    .Y(_02242_));
 sky130_fd_sc_hd__nand3_1 _08316_ (.A(_02240_),
    .B(_02143_),
    .C(_02242_),
    .Y(_02243_));
 sky130_fd_sc_hd__nand2_1 _08317_ (.A(_02230_),
    .B(\Qset[0][4] ),
    .Y(_02244_));
 sky130_fd_sc_hd__nand2_1 _08318_ (.A(_02141_),
    .B(\Qset[1][4] ),
    .Y(_02245_));
 sky130_fd_sc_hd__nand3_1 _08319_ (.A(_02244_),
    .B(_02147_),
    .C(_02245_),
    .Y(_02246_));
 sky130_fd_sc_hd__nand2_1 _08320_ (.A(_02243_),
    .B(_02246_),
    .Y(_02247_));
 sky130_fd_sc_hd__buf_4 _08321_ (.A(_02141_),
    .X(_02248_));
 sky130_fd_sc_hd__inv_2 _08322_ (.A(\Oset[2][4] ),
    .Y(_02249_));
 sky130_fd_sc_hd__clkbuf_4 _08323_ (.A(_02143_),
    .X(_02250_));
 sky130_fd_sc_hd__nand2_1 _08324_ (.A(_02248_),
    .B(\Oset[3][4] ),
    .Y(_02251_));
 sky130_fd_sc_hd__o211ai_1 _08325_ (.A1(_02248_),
    .A2(_02249_),
    .B1(_02250_),
    .C1(_02251_),
    .Y(_02252_));
 sky130_fd_sc_hd__inv_2 _08326_ (.A(\Oset[0][4] ),
    .Y(_02253_));
 sky130_fd_sc_hd__clkbuf_4 _08327_ (.A(_02147_),
    .X(_02254_));
 sky130_fd_sc_hd__nand2_1 _08328_ (.A(_02241_),
    .B(\Oset[1][4] ),
    .Y(_02255_));
 sky130_fd_sc_hd__o211ai_1 _08329_ (.A1(_02241_),
    .A2(_02253_),
    .B1(_02254_),
    .C1(_02255_),
    .Y(_02256_));
 sky130_fd_sc_hd__nand2_1 _08330_ (.A(_02252_),
    .B(_02256_),
    .Y(_02257_));
 sky130_fd_sc_hd__mux2_1 _08331_ (.A0(\H[2][4] ),
    .A1(\H[3][4] ),
    .S(_02241_),
    .X(_02258_));
 sky130_fd_sc_hd__nand2_1 _08332_ (.A(_02258_),
    .B(_02250_),
    .Y(_02259_));
 sky130_fd_sc_hd__buf_6 _08333_ (.A(_02230_),
    .X(_02260_));
 sky130_fd_sc_hd__buf_4 _08334_ (.A(_02141_),
    .X(_02261_));
 sky130_fd_sc_hd__o21a_1 _08335_ (.A1(_02261_),
    .A2(\H[0][4] ),
    .B1(_02254_),
    .X(_02262_));
 sky130_fd_sc_hd__o21ai_1 _08336_ (.A1(_02260_),
    .A2(\H[1][4] ),
    .B1(_02262_),
    .Y(_02263_));
 sky130_fd_sc_hd__a21o_2 _08337_ (.A1(_02259_),
    .A2(_02263_),
    .B1(_01552_),
    .X(_02264_));
 sky130_fd_sc_hd__o221ai_4 _08338_ (.A1(_02126_),
    .A2(_02247_),
    .B1(_02140_),
    .B2(_02257_),
    .C1(_02264_),
    .Y(_02265_));
 sky130_fd_sc_hd__mux2_1 _08339_ (.A0(_02265_),
    .A1(net58),
    .S(_02170_),
    .X(_02266_));
 sky130_fd_sc_hd__clkbuf_1 _08340_ (.A(_02266_),
    .X(_00232_));
 sky130_fd_sc_hd__nand2_1 _08341_ (.A(_02230_),
    .B(\Qset[2][5] ),
    .Y(_02267_));
 sky130_fd_sc_hd__nand2_1 _08342_ (.A(_02241_),
    .B(\Qset[3][5] ),
    .Y(_02268_));
 sky130_fd_sc_hd__nand3_1 _08343_ (.A(_02267_),
    .B(_02143_),
    .C(_02268_),
    .Y(_02269_));
 sky130_fd_sc_hd__nand2_1 _08344_ (.A(_02230_),
    .B(\Qset[0][5] ),
    .Y(_02270_));
 sky130_fd_sc_hd__nand2_1 _08345_ (.A(_02141_),
    .B(\Qset[1][5] ),
    .Y(_02271_));
 sky130_fd_sc_hd__nand3_1 _08346_ (.A(_02270_),
    .B(_02147_),
    .C(_02271_),
    .Y(_02272_));
 sky130_fd_sc_hd__nand2_1 _08347_ (.A(_02269_),
    .B(_02272_),
    .Y(_02273_));
 sky130_fd_sc_hd__inv_2 _08348_ (.A(\Oset[2][5] ),
    .Y(_02274_));
 sky130_fd_sc_hd__nor2_1 _08349_ (.A(_02241_),
    .B(_02274_),
    .Y(_02275_));
 sky130_fd_sc_hd__a211o_1 _08350_ (.A1(_02241_),
    .A2(\Oset[3][5] ),
    .B1(_02147_),
    .C1(_02275_),
    .X(_02276_));
 sky130_fd_sc_hd__inv_2 _08351_ (.A(\Oset[0][5] ),
    .Y(_02277_));
 sky130_fd_sc_hd__nor2_1 _08352_ (.A(_02141_),
    .B(_02277_),
    .Y(_02278_));
 sky130_fd_sc_hd__a211o_1 _08353_ (.A1(_02241_),
    .A2(\Oset[1][5] ),
    .B1(_02143_),
    .C1(_02278_),
    .X(_02279_));
 sky130_fd_sc_hd__nand2_1 _08354_ (.A(_02276_),
    .B(_02279_),
    .Y(_02280_));
 sky130_fd_sc_hd__inv_2 _08355_ (.A(\H[0][5] ),
    .Y(_02281_));
 sky130_fd_sc_hd__nor2_1 _08356_ (.A(\H[1][5] ),
    .B(_02230_),
    .Y(_02282_));
 sky130_fd_sc_hd__a211o_1 _08357_ (.A1(_02260_),
    .A2(_02281_),
    .B1(_02250_),
    .C1(_02282_),
    .X(_02283_));
 sky130_fd_sc_hd__o21a_1 _08358_ (.A1(_02261_),
    .A2(\H[2][5] ),
    .B1(_02250_),
    .X(_02284_));
 sky130_fd_sc_hd__o21ai_1 _08359_ (.A1(_02260_),
    .A2(\H[3][5] ),
    .B1(_02284_),
    .Y(_02285_));
 sky130_fd_sc_hd__a21o_2 _08360_ (.A1(_02283_),
    .A2(_02285_),
    .B1(_01552_),
    .X(_02286_));
 sky130_fd_sc_hd__o221ai_2 _08361_ (.A1(_02126_),
    .A2(_02273_),
    .B1(_02140_),
    .B2(_02280_),
    .C1(_02286_),
    .Y(_02287_));
 sky130_fd_sc_hd__mux2_1 _08362_ (.A0(_02287_),
    .A1(net59),
    .S(_02170_),
    .X(_02288_));
 sky130_fd_sc_hd__clkbuf_1 _08363_ (.A(_02288_),
    .X(_00233_));
 sky130_fd_sc_hd__inv_2 _08364_ (.A(\Qset[2][6] ),
    .Y(_02289_));
 sky130_fd_sc_hd__nand2_1 _08365_ (.A(_02261_),
    .B(\Qset[3][6] ),
    .Y(_02290_));
 sky130_fd_sc_hd__o211ai_1 _08366_ (.A1(_02248_),
    .A2(_02289_),
    .B1(_02250_),
    .C1(_02290_),
    .Y(_02291_));
 sky130_fd_sc_hd__inv_2 _08367_ (.A(\Qset[0][6] ),
    .Y(_02292_));
 sky130_fd_sc_hd__nand2_1 _08368_ (.A(_02248_),
    .B(\Qset[1][6] ),
    .Y(_02293_));
 sky130_fd_sc_hd__o211ai_1 _08369_ (.A1(_02248_),
    .A2(_02292_),
    .B1(_02254_),
    .C1(_02293_),
    .Y(_02294_));
 sky130_fd_sc_hd__nand2_2 _08370_ (.A(_02291_),
    .B(_02294_),
    .Y(_02295_));
 sky130_fd_sc_hd__inv_2 _08371_ (.A(\Oset[2][6] ),
    .Y(_02296_));
 sky130_fd_sc_hd__nor2_1 _08372_ (.A(_02248_),
    .B(_02296_),
    .Y(_02297_));
 sky130_fd_sc_hd__a211o_1 _08373_ (.A1(_02261_),
    .A2(\Oset[3][6] ),
    .B1(_02254_),
    .C1(_02297_),
    .X(_02298_));
 sky130_fd_sc_hd__inv_2 _08374_ (.A(\Oset[0][6] ),
    .Y(_02299_));
 sky130_fd_sc_hd__nor2_1 _08375_ (.A(_02248_),
    .B(_02299_),
    .Y(_02300_));
 sky130_fd_sc_hd__a211o_1 _08376_ (.A1(_02261_),
    .A2(\Oset[1][6] ),
    .B1(_02250_),
    .C1(_02300_),
    .X(_02301_));
 sky130_fd_sc_hd__nand2_2 _08377_ (.A(_02298_),
    .B(_02301_),
    .Y(_02302_));
 sky130_fd_sc_hd__inv_2 _08378_ (.A(\H[0][6] ),
    .Y(_02303_));
 sky130_fd_sc_hd__nor2_1 _08379_ (.A(\H[1][6] ),
    .B(_02260_),
    .Y(_02304_));
 sky130_fd_sc_hd__a211o_1 _08380_ (.A1(_02260_),
    .A2(_02303_),
    .B1(_02250_),
    .C1(_02304_),
    .X(_02305_));
 sky130_fd_sc_hd__o21a_1 _08381_ (.A1(_02261_),
    .A2(\H[2][6] ),
    .B1(_02250_),
    .X(_02306_));
 sky130_fd_sc_hd__o21ai_1 _08382_ (.A1(_02260_),
    .A2(\H[3][6] ),
    .B1(_02306_),
    .Y(_02307_));
 sky130_fd_sc_hd__a21o_2 _08383_ (.A1(_02305_),
    .A2(_02307_),
    .B1(_01552_),
    .X(_02308_));
 sky130_fd_sc_hd__o221ai_4 _08384_ (.A1(_02126_),
    .A2(_02295_),
    .B1(_02140_),
    .B2(_02302_),
    .C1(_02308_),
    .Y(_02309_));
 sky130_fd_sc_hd__mux2_1 _08385_ (.A0(_02309_),
    .A1(net60),
    .S(_02170_),
    .X(_02310_));
 sky130_fd_sc_hd__clkbuf_1 _08386_ (.A(_02310_),
    .X(_00234_));
 sky130_fd_sc_hd__buf_8 _08387_ (.A(_00591_),
    .X(_02311_));
 sky130_fd_sc_hd__inv_2 _08388_ (.A(\Qset[2][7] ),
    .Y(_02312_));
 sky130_fd_sc_hd__nor2_1 _08389_ (.A(_02241_),
    .B(_02312_),
    .Y(_02313_));
 sky130_fd_sc_hd__a211o_1 _08390_ (.A1(_02248_),
    .A2(\Qset[3][7] ),
    .B1(_02254_),
    .C1(_02313_),
    .X(_02314_));
 sky130_fd_sc_hd__inv_2 _08391_ (.A(\Qset[0][7] ),
    .Y(_02315_));
 sky130_fd_sc_hd__nor2_1 _08392_ (.A(_02241_),
    .B(_02315_),
    .Y(_02316_));
 sky130_fd_sc_hd__a211o_1 _08393_ (.A1(_02248_),
    .A2(\Qset[1][7] ),
    .B1(_02143_),
    .C1(_02316_),
    .X(_02317_));
 sky130_fd_sc_hd__nand2_2 _08394_ (.A(_02314_),
    .B(_02317_),
    .Y(_02318_));
 sky130_fd_sc_hd__buf_4 _08395_ (.A(_02248_),
    .X(_02319_));
 sky130_fd_sc_hd__inv_2 _08396_ (.A(\Oset[2][7] ),
    .Y(_02320_));
 sky130_fd_sc_hd__nor2_1 _08397_ (.A(_02261_),
    .B(_02320_),
    .Y(_02321_));
 sky130_fd_sc_hd__a211o_1 _08398_ (.A1(_02319_),
    .A2(\Oset[3][7] ),
    .B1(_02254_),
    .C1(_02321_),
    .X(_02322_));
 sky130_fd_sc_hd__inv_2 _08399_ (.A(\Oset[0][7] ),
    .Y(_02323_));
 sky130_fd_sc_hd__nor2_1 _08400_ (.A(_02261_),
    .B(_02323_),
    .Y(_02324_));
 sky130_fd_sc_hd__a211o_1 _08401_ (.A1(_02319_),
    .A2(\Oset[1][7] ),
    .B1(_02250_),
    .C1(_02324_),
    .X(_02325_));
 sky130_fd_sc_hd__nand2_2 _08402_ (.A(_02322_),
    .B(_02325_),
    .Y(_02326_));
 sky130_fd_sc_hd__clkbuf_4 _08403_ (.A(_02260_),
    .X(_02327_));
 sky130_fd_sc_hd__buf_4 _08404_ (.A(_02261_),
    .X(_02328_));
 sky130_fd_sc_hd__clkbuf_4 _08405_ (.A(_02250_),
    .X(_02329_));
 sky130_fd_sc_hd__o21a_1 _08406_ (.A1(_02328_),
    .A2(\H[2][7] ),
    .B1(_02329_),
    .X(_02330_));
 sky130_fd_sc_hd__o21ai_1 _08407_ (.A1(_02327_),
    .A2(\H[3][7] ),
    .B1(_02330_),
    .Y(_02331_));
 sky130_fd_sc_hd__o21a_1 _08408_ (.A1(_02319_),
    .A2(\H[0][7] ),
    .B1(_02254_),
    .X(_02332_));
 sky130_fd_sc_hd__o21ai_1 _08409_ (.A1(_02327_),
    .A2(\H[1][7] ),
    .B1(_02332_),
    .Y(_02333_));
 sky130_fd_sc_hd__a21o_2 _08410_ (.A1(_02331_),
    .A2(_02333_),
    .B1(_01552_),
    .X(_02334_));
 sky130_fd_sc_hd__o221ai_4 _08411_ (.A1(_02311_),
    .A2(_02318_),
    .B1(_02140_),
    .B2(_02326_),
    .C1(_02334_),
    .Y(_02335_));
 sky130_fd_sc_hd__mux2_1 _08412_ (.A0(_02335_),
    .A1(net61),
    .S(_02170_),
    .X(_02336_));
 sky130_fd_sc_hd__clkbuf_1 _08413_ (.A(_02336_),
    .X(_00235_));
 sky130_fd_sc_hd__nor2_1 _08414_ (.A(\Qset[3][8] ),
    .B(_02260_),
    .Y(_02337_));
 sky130_fd_sc_hd__o21ai_1 _08415_ (.A1(_02319_),
    .A2(\Qset[2][8] ),
    .B1(_02329_),
    .Y(_02338_));
 sky130_fd_sc_hd__nor2_1 _08416_ (.A(_02319_),
    .B(\Qset[0][8] ),
    .Y(_02339_));
 sky130_fd_sc_hd__o21ai_1 _08417_ (.A1(\Qset[1][8] ),
    .A2(_02260_),
    .B1(_02254_),
    .Y(_02340_));
 sky130_fd_sc_hd__o22a_2 _08418_ (.A1(_02337_),
    .A2(_02338_),
    .B1(_02339_),
    .B2(_02340_),
    .X(_02341_));
 sky130_fd_sc_hd__mux2_1 _08419_ (.A0(\Oset[2][8] ),
    .A1(\Oset[3][8] ),
    .S(_02261_),
    .X(_02342_));
 sky130_fd_sc_hd__nor2_1 _08420_ (.A(_02319_),
    .B(\Oset[0][8] ),
    .Y(_02343_));
 sky130_fd_sc_hd__o21ai_1 _08421_ (.A1(\Oset[1][8] ),
    .A2(_02260_),
    .B1(_02254_),
    .Y(_02344_));
 sky130_fd_sc_hd__o2bb2a_2 _08422_ (.A1_N(_02329_),
    .A2_N(_02342_),
    .B1(_02343_),
    .B2(_02344_),
    .X(_02345_));
 sky130_fd_sc_hd__inv_2 _08423_ (.A(\H[2][8] ),
    .Y(_02346_));
 sky130_fd_sc_hd__clkbuf_4 _08424_ (.A(_02254_),
    .X(_02347_));
 sky130_fd_sc_hd__nor2_1 _08425_ (.A(\H[3][8] ),
    .B(_02327_),
    .Y(_02348_));
 sky130_fd_sc_hd__a211o_1 _08426_ (.A1(_02327_),
    .A2(_02346_),
    .B1(_02347_),
    .C1(_02348_),
    .X(_02349_));
 sky130_fd_sc_hd__inv_2 _08427_ (.A(\H[0][8] ),
    .Y(_02350_));
 sky130_fd_sc_hd__nor2_1 _08428_ (.A(\H[1][8] ),
    .B(_02327_),
    .Y(_02351_));
 sky130_fd_sc_hd__a211o_1 _08429_ (.A1(_02327_),
    .A2(_02350_),
    .B1(_02329_),
    .C1(_02351_),
    .X(_02352_));
 sky130_fd_sc_hd__a21o_1 _08430_ (.A1(_02349_),
    .A2(_02352_),
    .B1(_01553_),
    .X(_02353_));
 sky130_fd_sc_hd__o221ai_4 _08431_ (.A1(_02311_),
    .A2(_02341_),
    .B1(_02140_),
    .B2(_02345_),
    .C1(_02353_),
    .Y(_02354_));
 sky130_fd_sc_hd__mux2_1 _08432_ (.A0(_02354_),
    .A1(net62),
    .S(_02170_),
    .X(_02355_));
 sky130_fd_sc_hd__clkbuf_1 _08433_ (.A(_02355_),
    .X(_00236_));
 sky130_fd_sc_hd__buf_4 _08434_ (.A(_02319_),
    .X(_02356_));
 sky130_fd_sc_hd__inv_2 _08435_ (.A(\Qset[2][9] ),
    .Y(_02357_));
 sky130_fd_sc_hd__nor2_1 _08436_ (.A(_02328_),
    .B(_02357_),
    .Y(_02358_));
 sky130_fd_sc_hd__a211o_1 _08437_ (.A1(_02356_),
    .A2(\Qset[3][9] ),
    .B1(_02347_),
    .C1(_02358_),
    .X(_02359_));
 sky130_fd_sc_hd__inv_2 _08438_ (.A(\Qset[0][9] ),
    .Y(_02360_));
 sky130_fd_sc_hd__nor2_1 _08439_ (.A(_02328_),
    .B(_02360_),
    .Y(_02361_));
 sky130_fd_sc_hd__a211o_1 _08440_ (.A1(_02356_),
    .A2(\Qset[1][9] ),
    .B1(_02329_),
    .C1(_02361_),
    .X(_02362_));
 sky130_fd_sc_hd__nand2_2 _08441_ (.A(_02359_),
    .B(_02362_),
    .Y(_02363_));
 sky130_fd_sc_hd__buf_4 _08442_ (.A(_02328_),
    .X(_02364_));
 sky130_fd_sc_hd__inv_2 _08443_ (.A(\Oset[2][9] ),
    .Y(_02365_));
 sky130_fd_sc_hd__nor2_1 _08444_ (.A(_02356_),
    .B(_02365_),
    .Y(_02366_));
 sky130_fd_sc_hd__a211o_1 _08445_ (.A1(_02364_),
    .A2(\Oset[3][9] ),
    .B1(_02347_),
    .C1(_02366_),
    .X(_02367_));
 sky130_fd_sc_hd__inv_2 _08446_ (.A(\Oset[0][9] ),
    .Y(_02368_));
 sky130_fd_sc_hd__nor2_1 _08447_ (.A(_02356_),
    .B(_02368_),
    .Y(_02369_));
 sky130_fd_sc_hd__a211o_1 _08448_ (.A1(_02356_),
    .A2(\Oset[1][9] ),
    .B1(_02329_),
    .C1(_02369_),
    .X(_02370_));
 sky130_fd_sc_hd__nand2_2 _08449_ (.A(_02367_),
    .B(_02370_),
    .Y(_02371_));
 sky130_fd_sc_hd__inv_2 _08450_ (.A(\H[3][9] ),
    .Y(_02372_));
 sky130_fd_sc_hd__buf_4 _08451_ (.A(_02364_),
    .X(_02373_));
 sky130_fd_sc_hd__clkbuf_4 _08452_ (.A(_02347_),
    .X(_02374_));
 sky130_fd_sc_hd__nor2_1 _08453_ (.A(_02373_),
    .B(\H[2][9] ),
    .Y(_02375_));
 sky130_fd_sc_hd__a211o_1 _08454_ (.A1(_02372_),
    .A2(_02373_),
    .B1(_02374_),
    .C1(_02375_),
    .X(_02376_));
 sky130_fd_sc_hd__inv_2 _08455_ (.A(\H[1][9] ),
    .Y(_02377_));
 sky130_fd_sc_hd__buf_4 _08456_ (.A(_02329_),
    .X(_02378_));
 sky130_fd_sc_hd__nor2_1 _08457_ (.A(_02373_),
    .B(\H[0][9] ),
    .Y(_02379_));
 sky130_fd_sc_hd__a211o_1 _08458_ (.A1(_02377_),
    .A2(_02373_),
    .B1(_02378_),
    .C1(_02379_),
    .X(_02380_));
 sky130_fd_sc_hd__a21o_2 _08459_ (.A1(_02376_),
    .A2(_02380_),
    .B1(_01553_),
    .X(_02381_));
 sky130_fd_sc_hd__o221ai_4 _08460_ (.A1(_02311_),
    .A2(_02363_),
    .B1(_02140_),
    .B2(_02371_),
    .C1(_02381_),
    .Y(_02382_));
 sky130_fd_sc_hd__mux2_1 _08461_ (.A0(_02382_),
    .A1(net63),
    .S(_02170_),
    .X(_02383_));
 sky130_fd_sc_hd__clkbuf_1 _08462_ (.A(_02383_),
    .X(_00237_));
 sky130_fd_sc_hd__inv_2 _08463_ (.A(\Oset[2][10] ),
    .Y(_02384_));
 sky130_fd_sc_hd__nor2_1 _08464_ (.A(_02356_),
    .B(_02384_),
    .Y(_02385_));
 sky130_fd_sc_hd__a211o_1 _08465_ (.A1(_02364_),
    .A2(\Oset[3][10] ),
    .B1(_02347_),
    .C1(_02385_),
    .X(_02386_));
 sky130_fd_sc_hd__inv_2 _08466_ (.A(\Oset[0][10] ),
    .Y(_02387_));
 sky130_fd_sc_hd__nor2_1 _08467_ (.A(_02356_),
    .B(_02387_),
    .Y(_02388_));
 sky130_fd_sc_hd__a211o_1 _08468_ (.A1(_02364_),
    .A2(\Oset[1][10] ),
    .B1(_02378_),
    .C1(_02388_),
    .X(_02389_));
 sky130_fd_sc_hd__nand2_2 _08469_ (.A(_02386_),
    .B(_02389_),
    .Y(_02390_));
 sky130_fd_sc_hd__inv_2 _08470_ (.A(\Qset[0][10] ),
    .Y(_02391_));
 sky130_fd_sc_hd__nand2_1 _08471_ (.A(_02327_),
    .B(_02391_),
    .Y(_02392_));
 sky130_fd_sc_hd__o21a_1 _08472_ (.A1(\Qset[1][10] ),
    .A2(_02327_),
    .B1(_02347_),
    .X(_02393_));
 sky130_fd_sc_hd__mux2_1 _08473_ (.A0(\Qset[2][10] ),
    .A1(\Qset[3][10] ),
    .S(_02319_),
    .X(_02394_));
 sky130_fd_sc_hd__a22oi_4 _08474_ (.A1(_02392_),
    .A2(_02393_),
    .B1(_02394_),
    .B2(_02378_),
    .Y(_02395_));
 sky130_fd_sc_hd__inv_2 _08475_ (.A(\H[3][10] ),
    .Y(_02396_));
 sky130_fd_sc_hd__buf_4 _08476_ (.A(_02356_),
    .X(_02397_));
 sky130_fd_sc_hd__nor2_1 _08477_ (.A(_02397_),
    .B(\H[2][10] ),
    .Y(_02398_));
 sky130_fd_sc_hd__a211o_1 _08478_ (.A1(_02396_),
    .A2(_02373_),
    .B1(_02374_),
    .C1(_02398_),
    .X(_02399_));
 sky130_fd_sc_hd__inv_2 _08479_ (.A(\H[1][10] ),
    .Y(_02400_));
 sky130_fd_sc_hd__nor2_1 _08480_ (.A(_02397_),
    .B(\H[0][10] ),
    .Y(_02401_));
 sky130_fd_sc_hd__a211o_1 _08481_ (.A1(_02400_),
    .A2(_02397_),
    .B1(_02378_),
    .C1(_02401_),
    .X(_02402_));
 sky130_fd_sc_hd__a21o_2 _08482_ (.A1(_02399_),
    .A2(_02402_),
    .B1(_01553_),
    .X(_02403_));
 sky130_fd_sc_hd__o221ai_4 _08483_ (.A1(_02139_),
    .A2(_02390_),
    .B1(_02126_),
    .B2(_02395_),
    .C1(_02403_),
    .Y(_02404_));
 sky130_fd_sc_hd__mux2_1 _08484_ (.A0(_02404_),
    .A1(net49),
    .S(_02169_),
    .X(_02405_));
 sky130_fd_sc_hd__clkbuf_1 _08485_ (.A(_02405_),
    .X(_00238_));
 sky130_fd_sc_hd__inv_2 _08486_ (.A(\Qset[2][11] ),
    .Y(_02406_));
 sky130_fd_sc_hd__nor2_1 _08487_ (.A(_02328_),
    .B(_02406_),
    .Y(_02407_));
 sky130_fd_sc_hd__a211o_1 _08488_ (.A1(_02328_),
    .A2(\Qset[3][11] ),
    .B1(_02347_),
    .C1(_02407_),
    .X(_02408_));
 sky130_fd_sc_hd__inv_2 _08489_ (.A(\Qset[0][11] ),
    .Y(_02409_));
 sky130_fd_sc_hd__nor2_1 _08490_ (.A(_02319_),
    .B(_02409_),
    .Y(_02410_));
 sky130_fd_sc_hd__a211o_1 _08491_ (.A1(_02328_),
    .A2(\Qset[1][11] ),
    .B1(_02329_),
    .C1(_02410_),
    .X(_02411_));
 sky130_fd_sc_hd__nand2_2 _08492_ (.A(_02408_),
    .B(_02411_),
    .Y(_02412_));
 sky130_fd_sc_hd__inv_2 _08493_ (.A(\Oset[2][11] ),
    .Y(_02413_));
 sky130_fd_sc_hd__nor2_1 _08494_ (.A(_02356_),
    .B(_02413_),
    .Y(_02414_));
 sky130_fd_sc_hd__a211o_1 _08495_ (.A1(_02364_),
    .A2(\Oset[3][11] ),
    .B1(_02347_),
    .C1(_02414_),
    .X(_02415_));
 sky130_fd_sc_hd__inv_2 _08496_ (.A(\Oset[0][11] ),
    .Y(_02416_));
 sky130_fd_sc_hd__nor2_1 _08497_ (.A(_02356_),
    .B(_02416_),
    .Y(_02417_));
 sky130_fd_sc_hd__a211o_1 _08498_ (.A1(_02364_),
    .A2(\Oset[1][11] ),
    .B1(_02329_),
    .C1(_02417_),
    .X(_02418_));
 sky130_fd_sc_hd__nand2_2 _08499_ (.A(_02415_),
    .B(_02418_),
    .Y(_02419_));
 sky130_fd_sc_hd__inv_2 _08500_ (.A(\H[3][11] ),
    .Y(_02420_));
 sky130_fd_sc_hd__nor2_1 _08501_ (.A(_02397_),
    .B(\H[2][11] ),
    .Y(_02421_));
 sky130_fd_sc_hd__a211o_1 _08502_ (.A1(_02420_),
    .A2(_02373_),
    .B1(_02374_),
    .C1(_02421_),
    .X(_02422_));
 sky130_fd_sc_hd__inv_2 _08503_ (.A(\H[1][11] ),
    .Y(_02423_));
 sky130_fd_sc_hd__nor2_1 _08504_ (.A(_02397_),
    .B(\H[0][11] ),
    .Y(_02424_));
 sky130_fd_sc_hd__a211o_1 _08505_ (.A1(_02423_),
    .A2(_02373_),
    .B1(_02378_),
    .C1(_02424_),
    .X(_02425_));
 sky130_fd_sc_hd__a21o_2 _08506_ (.A1(_02422_),
    .A2(_02425_),
    .B1(_01553_),
    .X(_02426_));
 sky130_fd_sc_hd__o221ai_4 _08507_ (.A1(_02311_),
    .A2(_02412_),
    .B1(_02139_),
    .B2(_02419_),
    .C1(_02426_),
    .Y(_02427_));
 sky130_fd_sc_hd__mux2_1 _08508_ (.A0(_02427_),
    .A1(net50),
    .S(_02169_),
    .X(_02428_));
 sky130_fd_sc_hd__clkbuf_1 _08509_ (.A(_02428_),
    .X(_00239_));
 sky130_fd_sc_hd__inv_2 _08510_ (.A(\Qset[2][12] ),
    .Y(_02429_));
 sky130_fd_sc_hd__nor2_1 _08511_ (.A(_02328_),
    .B(_02429_),
    .Y(_02430_));
 sky130_fd_sc_hd__a211o_1 _08512_ (.A1(_02328_),
    .A2(\Qset[3][12] ),
    .B1(_02347_),
    .C1(_02430_),
    .X(_02431_));
 sky130_fd_sc_hd__inv_2 _08513_ (.A(\Qset[0][12] ),
    .Y(_02432_));
 sky130_fd_sc_hd__nor2_1 _08514_ (.A(_02319_),
    .B(_02432_),
    .Y(_02433_));
 sky130_fd_sc_hd__a211o_1 _08515_ (.A1(_02328_),
    .A2(\Qset[1][12] ),
    .B1(_02329_),
    .C1(_02433_),
    .X(_02434_));
 sky130_fd_sc_hd__nand2_2 _08516_ (.A(_02431_),
    .B(_02434_),
    .Y(_02435_));
 sky130_fd_sc_hd__inv_2 _08517_ (.A(\Oset[2][12] ),
    .Y(_02436_));
 sky130_fd_sc_hd__nor2_1 _08518_ (.A(_02364_),
    .B(_02436_),
    .Y(_02437_));
 sky130_fd_sc_hd__a211o_1 _08519_ (.A1(_02364_),
    .A2(\Oset[3][12] ),
    .B1(_02347_),
    .C1(_02437_),
    .X(_02438_));
 sky130_fd_sc_hd__inv_2 _08520_ (.A(\Oset[0][12] ),
    .Y(_02439_));
 sky130_fd_sc_hd__nor2_1 _08521_ (.A(_02364_),
    .B(_02439_),
    .Y(_02440_));
 sky130_fd_sc_hd__a211o_1 _08522_ (.A1(_02364_),
    .A2(\Oset[1][12] ),
    .B1(_02378_),
    .C1(_02440_),
    .X(_02441_));
 sky130_fd_sc_hd__nand2_1 _08523_ (.A(_02438_),
    .B(_02441_),
    .Y(_02442_));
 sky130_fd_sc_hd__mux2_1 _08524_ (.A0(\H[2][12] ),
    .A1(\H[3][12] ),
    .S(_02397_),
    .X(_02443_));
 sky130_fd_sc_hd__clkbuf_4 _08525_ (.A(_02378_),
    .X(_02444_));
 sky130_fd_sc_hd__nand2_1 _08526_ (.A(_02443_),
    .B(_02444_),
    .Y(_02445_));
 sky130_fd_sc_hd__inv_2 _08527_ (.A(\H[1][12] ),
    .Y(_02446_));
 sky130_fd_sc_hd__nor2_1 _08528_ (.A(_02373_),
    .B(\H[0][12] ),
    .Y(_02447_));
 sky130_fd_sc_hd__a211o_1 _08529_ (.A1(_02446_),
    .A2(_02373_),
    .B1(_02378_),
    .C1(_02447_),
    .X(_02448_));
 sky130_fd_sc_hd__a21o_2 _08530_ (.A1(_02445_),
    .A2(_02448_),
    .B1(_01553_),
    .X(_02449_));
 sky130_fd_sc_hd__o221ai_4 _08531_ (.A1(_02311_),
    .A2(_02435_),
    .B1(_02139_),
    .B2(_02442_),
    .C1(_02449_),
    .Y(_02450_));
 sky130_fd_sc_hd__mux2_1 _08532_ (.A0(_02450_),
    .A1(net51),
    .S(_02169_),
    .X(_02451_));
 sky130_fd_sc_hd__clkbuf_1 _08533_ (.A(_02451_),
    .X(_00240_));
 sky130_fd_sc_hd__inv_2 _08534_ (.A(\Qset[2][13] ),
    .Y(_02452_));
 sky130_fd_sc_hd__nor2_1 _08535_ (.A(_02397_),
    .B(_02452_),
    .Y(_02453_));
 sky130_fd_sc_hd__a211o_1 _08536_ (.A1(_02397_),
    .A2(\Qset[3][13] ),
    .B1(_02374_),
    .C1(_02453_),
    .X(_02454_));
 sky130_fd_sc_hd__inv_2 _08537_ (.A(\Qset[0][13] ),
    .Y(_02455_));
 sky130_fd_sc_hd__nor2_1 _08538_ (.A(_02397_),
    .B(_02455_),
    .Y(_02456_));
 sky130_fd_sc_hd__a211o_1 _08539_ (.A1(_02397_),
    .A2(\Qset[1][13] ),
    .B1(_02378_),
    .C1(_02456_),
    .X(_02457_));
 sky130_fd_sc_hd__nand2_1 _08540_ (.A(_02454_),
    .B(_02457_),
    .Y(_02458_));
 sky130_fd_sc_hd__buf_4 _08541_ (.A(_02373_),
    .X(_02459_));
 sky130_fd_sc_hd__inv_2 _08542_ (.A(\Oset[2][13] ),
    .Y(_02460_));
 sky130_fd_sc_hd__nor2_1 _08543_ (.A(_02459_),
    .B(_02460_),
    .Y(_02461_));
 sky130_fd_sc_hd__a211o_1 _08544_ (.A1(_02459_),
    .A2(\Oset[3][13] ),
    .B1(_02374_),
    .C1(_02461_),
    .X(_02462_));
 sky130_fd_sc_hd__inv_2 _08545_ (.A(\Oset[0][13] ),
    .Y(_02463_));
 sky130_fd_sc_hd__nor2_1 _08546_ (.A(_02459_),
    .B(_02463_),
    .Y(_02464_));
 sky130_fd_sc_hd__a211o_1 _08547_ (.A1(_02459_),
    .A2(\Oset[1][13] ),
    .B1(_02378_),
    .C1(_02464_),
    .X(_02465_));
 sky130_fd_sc_hd__nand2_1 _08548_ (.A(_02462_),
    .B(_02465_),
    .Y(_02466_));
 sky130_fd_sc_hd__mux2_1 _08549_ (.A0(\H[2][13] ),
    .A1(\H[3][13] ),
    .S(_02459_),
    .X(_02467_));
 sky130_fd_sc_hd__nand2_1 _08550_ (.A(_02467_),
    .B(_02444_),
    .Y(_02468_));
 sky130_fd_sc_hd__inv_2 _08551_ (.A(\H[1][13] ),
    .Y(_02469_));
 sky130_fd_sc_hd__buf_4 _08552_ (.A(_02459_),
    .X(_02470_));
 sky130_fd_sc_hd__nor2_1 _08553_ (.A(_02470_),
    .B(\H[0][13] ),
    .Y(_02471_));
 sky130_fd_sc_hd__a211o_1 _08554_ (.A1(_02469_),
    .A2(_02470_),
    .B1(_02444_),
    .C1(_02471_),
    .X(_02472_));
 sky130_fd_sc_hd__a21o_1 _08555_ (.A1(_02468_),
    .A2(_02472_),
    .B1(_01554_),
    .X(_02473_));
 sky130_fd_sc_hd__o221ai_4 _08556_ (.A1(_02311_),
    .A2(_02458_),
    .B1(_02139_),
    .B2(_02466_),
    .C1(_02473_),
    .Y(_02474_));
 sky130_fd_sc_hd__mux2_1 _08557_ (.A0(_02474_),
    .A1(net52),
    .S(_02169_),
    .X(_02475_));
 sky130_fd_sc_hd__clkbuf_1 _08558_ (.A(_02475_),
    .X(_00241_));
 sky130_fd_sc_hd__inv_2 _08559_ (.A(\Qset[2][14] ),
    .Y(_02476_));
 sky130_fd_sc_hd__nor2_1 _08560_ (.A(_02459_),
    .B(_02476_),
    .Y(_02477_));
 sky130_fd_sc_hd__a211o_1 _08561_ (.A1(_02459_),
    .A2(\Qset[3][14] ),
    .B1(_02374_),
    .C1(_02477_),
    .X(_02478_));
 sky130_fd_sc_hd__inv_2 _08562_ (.A(\Qset[0][14] ),
    .Y(_02479_));
 sky130_fd_sc_hd__nor2_1 _08563_ (.A(_02459_),
    .B(_02479_),
    .Y(_02480_));
 sky130_fd_sc_hd__a211o_1 _08564_ (.A1(_02459_),
    .A2(\Qset[1][14] ),
    .B1(_02444_),
    .C1(_02480_),
    .X(_02481_));
 sky130_fd_sc_hd__nand2_2 _08565_ (.A(_02478_),
    .B(_02481_),
    .Y(_02482_));
 sky130_fd_sc_hd__inv_2 _08566_ (.A(\Oset[2][14] ),
    .Y(_02483_));
 sky130_fd_sc_hd__nor2_1 _08567_ (.A(_02470_),
    .B(_02483_),
    .Y(_02484_));
 sky130_fd_sc_hd__a211o_1 _08568_ (.A1(_02470_),
    .A2(\Oset[3][14] ),
    .B1(_02374_),
    .C1(_02484_),
    .X(_02485_));
 sky130_fd_sc_hd__inv_2 _08569_ (.A(\Oset[0][14] ),
    .Y(_02486_));
 sky130_fd_sc_hd__nor2_1 _08570_ (.A(_02470_),
    .B(_02486_),
    .Y(_02487_));
 sky130_fd_sc_hd__a211o_1 _08571_ (.A1(_02470_),
    .A2(\Oset[1][14] ),
    .B1(_02444_),
    .C1(_02487_),
    .X(_02488_));
 sky130_fd_sc_hd__nand2_1 _08572_ (.A(_02485_),
    .B(_02488_),
    .Y(_02489_));
 sky130_fd_sc_hd__inv_2 _08573_ (.A(\H[3][14] ),
    .Y(_02490_));
 sky130_fd_sc_hd__buf_4 _08574_ (.A(_02470_),
    .X(_02491_));
 sky130_fd_sc_hd__nor2_1 _08575_ (.A(_02491_),
    .B(\H[2][14] ),
    .Y(_02492_));
 sky130_fd_sc_hd__a211o_1 _08576_ (.A1(_02490_),
    .A2(_02491_),
    .B1(_02374_),
    .C1(_02492_),
    .X(_02493_));
 sky130_fd_sc_hd__inv_2 _08577_ (.A(\H[1][14] ),
    .Y(_02494_));
 sky130_fd_sc_hd__nor2_1 _08578_ (.A(_02470_),
    .B(\H[0][14] ),
    .Y(_02495_));
 sky130_fd_sc_hd__a211o_1 _08579_ (.A1(_02494_),
    .A2(_02491_),
    .B1(_02444_),
    .C1(_02495_),
    .X(_02496_));
 sky130_fd_sc_hd__a21o_2 _08580_ (.A1(_02493_),
    .A2(_02496_),
    .B1(_01554_),
    .X(_02497_));
 sky130_fd_sc_hd__o221ai_4 _08581_ (.A1(_02311_),
    .A2(_02482_),
    .B1(_02139_),
    .B2(_02489_),
    .C1(_02497_),
    .Y(_02498_));
 sky130_fd_sc_hd__mux2_1 _08582_ (.A0(_02498_),
    .A1(net53),
    .S(_02169_),
    .X(_02499_));
 sky130_fd_sc_hd__clkbuf_1 _08583_ (.A(_02499_),
    .X(_00242_));
 sky130_fd_sc_hd__inv_2 _08584_ (.A(\Qset[2][15] ),
    .Y(_02500_));
 sky130_fd_sc_hd__nor2_1 _08585_ (.A(_02470_),
    .B(_02500_),
    .Y(_02501_));
 sky130_fd_sc_hd__a211o_1 _08586_ (.A1(_02491_),
    .A2(\Qset[3][15] ),
    .B1(_02374_),
    .C1(_02501_),
    .X(_02502_));
 sky130_fd_sc_hd__inv_2 _08587_ (.A(\Qset[0][15] ),
    .Y(_02503_));
 sky130_fd_sc_hd__nor2_1 _08588_ (.A(_02470_),
    .B(_02503_),
    .Y(_02504_));
 sky130_fd_sc_hd__a211o_1 _08589_ (.A1(_02491_),
    .A2(\Qset[1][15] ),
    .B1(_02444_),
    .C1(_02504_),
    .X(_02505_));
 sky130_fd_sc_hd__nand2_2 _08590_ (.A(_02502_),
    .B(_02505_),
    .Y(_02506_));
 sky130_fd_sc_hd__inv_2 _08591_ (.A(\Oset[2][15] ),
    .Y(_02507_));
 sky130_fd_sc_hd__nor2_1 _08592_ (.A(_02491_),
    .B(_02507_),
    .Y(_02508_));
 sky130_fd_sc_hd__a211o_1 _08593_ (.A1(_02491_),
    .A2(\Oset[3][15] ),
    .B1(_02374_),
    .C1(_02508_),
    .X(_02509_));
 sky130_fd_sc_hd__inv_2 _08594_ (.A(\Oset[0][15] ),
    .Y(_02510_));
 sky130_fd_sc_hd__nor2_1 _08595_ (.A(_02491_),
    .B(_02510_),
    .Y(_02511_));
 sky130_fd_sc_hd__a211o_1 _08596_ (.A1(_02491_),
    .A2(\Oset[1][15] ),
    .B1(_02444_),
    .C1(_02511_),
    .X(_02512_));
 sky130_fd_sc_hd__nand2_1 _08597_ (.A(_02509_),
    .B(_02512_),
    .Y(_02513_));
 sky130_fd_sc_hd__inv_2 _08598_ (.A(\H[0][15] ),
    .Y(_02514_));
 sky130_fd_sc_hd__nor2_1 _08599_ (.A(\H[1][15] ),
    .B(_02327_),
    .Y(_02515_));
 sky130_fd_sc_hd__a211o_1 _08600_ (.A1(_02327_),
    .A2(_02514_),
    .B1(_02444_),
    .C1(_02515_),
    .X(_02516_));
 sky130_fd_sc_hd__mux2_1 _08601_ (.A0(\H[2][15] ),
    .A1(\H[3][15] ),
    .S(_02491_),
    .X(_02517_));
 sky130_fd_sc_hd__nand2_1 _08602_ (.A(_02517_),
    .B(_02444_),
    .Y(_02518_));
 sky130_fd_sc_hd__a21o_1 _08603_ (.A1(_02516_),
    .A2(_02518_),
    .B1(_01554_),
    .X(_02519_));
 sky130_fd_sc_hd__o221ai_4 _08604_ (.A1(_02311_),
    .A2(_02506_),
    .B1(_02139_),
    .B2(_02513_),
    .C1(_02519_),
    .Y(_02520_));
 sky130_fd_sc_hd__mux2_1 _08605_ (.A0(_02520_),
    .A1(net54),
    .S(_02169_),
    .X(_02521_));
 sky130_fd_sc_hd__clkbuf_1 _08606_ (.A(_02521_),
    .X(_00243_));
 sky130_fd_sc_hd__clkinv_4 _08607_ (.A(_00006_),
    .Y(_02522_));
 sky130_fd_sc_hd__buf_4 _08608_ (.A(_02522_),
    .X(_02523_));
 sky130_fd_sc_hd__nand2_1 _08609_ (.A(_02523_),
    .B(\Qset[2][0] ),
    .Y(_02524_));
 sky130_fd_sc_hd__clkbuf_8 _08610_ (.A(_00007_),
    .X(_02525_));
 sky130_fd_sc_hd__clkbuf_8 _08611_ (.A(_02525_),
    .X(_02526_));
 sky130_fd_sc_hd__buf_6 _08612_ (.A(_00006_),
    .X(_02527_));
 sky130_fd_sc_hd__buf_6 _08613_ (.A(_02527_),
    .X(_02528_));
 sky130_fd_sc_hd__buf_6 _08614_ (.A(_02528_),
    .X(_02529_));
 sky130_fd_sc_hd__nand2_1 _08615_ (.A(\Qset[3][0] ),
    .B(_02529_),
    .Y(_02530_));
 sky130_fd_sc_hd__nand3_1 _08616_ (.A(_02524_),
    .B(_02526_),
    .C(_02530_),
    .Y(_02531_));
 sky130_fd_sc_hd__nand2_1 _08617_ (.A(_02523_),
    .B(\Qset[0][0] ),
    .Y(_02532_));
 sky130_fd_sc_hd__inv_2 _08618_ (.A(_00007_),
    .Y(_02533_));
 sky130_fd_sc_hd__buf_6 _08619_ (.A(_02533_),
    .X(_02534_));
 sky130_fd_sc_hd__clkbuf_8 _08620_ (.A(_02534_),
    .X(_02535_));
 sky130_fd_sc_hd__nand2_1 _08621_ (.A(\Qset[1][0] ),
    .B(_02529_),
    .Y(_02536_));
 sky130_fd_sc_hd__nand3_1 _08622_ (.A(_02532_),
    .B(_02535_),
    .C(_02536_),
    .Y(_02537_));
 sky130_fd_sc_hd__nand2_1 _08623_ (.A(_02531_),
    .B(_02537_),
    .Y(_02538_));
 sky130_fd_sc_hd__nor2_4 _08624_ (.A(Oreg3),
    .B(Oreg2),
    .Y(_02539_));
 sky130_fd_sc_hd__buf_4 _08625_ (.A(_02539_),
    .X(_02540_));
 sky130_fd_sc_hd__o21ai_1 _08626_ (.A1(_01959_),
    .A2(_00580_),
    .B1(_02540_),
    .Y(_02541_));
 sky130_fd_sc_hd__inv_2 _08627_ (.A(_02541_),
    .Y(_02542_));
 sky130_fd_sc_hd__o21ai_1 _08628_ (.A1(_02161_),
    .A2(_02538_),
    .B1(_02542_),
    .Y(_02543_));
 sky130_fd_sc_hd__buf_6 _08629_ (.A(_02527_),
    .X(_02544_));
 sky130_fd_sc_hd__buf_4 _08630_ (.A(_02544_),
    .X(_02545_));
 sky130_fd_sc_hd__nand2_1 _08631_ (.A(\Oset[3][0] ),
    .B(_02545_),
    .Y(_02546_));
 sky130_fd_sc_hd__o211ai_1 _08632_ (.A1(_02545_),
    .A2(_02142_),
    .B1(_02526_),
    .C1(_02546_),
    .Y(_02547_));
 sky130_fd_sc_hd__nand2_1 _08633_ (.A(\Oset[1][0] ),
    .B(_02529_),
    .Y(_02548_));
 sky130_fd_sc_hd__o211ai_1 _08634_ (.A1(_02545_),
    .A2(_02146_),
    .B1(_02535_),
    .C1(_02548_),
    .Y(_02549_));
 sky130_fd_sc_hd__nand2_2 _08635_ (.A(_02547_),
    .B(_02549_),
    .Y(_02550_));
 sky130_fd_sc_hd__inv_2 _08636_ (.A(_02539_),
    .Y(_02551_));
 sky130_fd_sc_hd__buf_2 _08637_ (.A(_02551_),
    .X(_02552_));
 sky130_fd_sc_hd__nand2_1 _08638_ (.A(_02550_),
    .B(_02552_),
    .Y(_02553_));
 sky130_fd_sc_hd__nand2_1 _08639_ (.A(_02543_),
    .B(_02553_),
    .Y(_02554_));
 sky130_fd_sc_hd__nor2_4 _08640_ (.A(Hreg3),
    .B(Hreg2),
    .Y(_02555_));
 sky130_fd_sc_hd__buf_4 _08641_ (.A(_02555_),
    .X(_02556_));
 sky130_fd_sc_hd__o21ai_1 _08642_ (.A1(_01959_),
    .A2(_01154_),
    .B1(_02556_),
    .Y(_02557_));
 sky130_fd_sc_hd__inv_2 _08643_ (.A(_02557_),
    .Y(_02558_));
 sky130_fd_sc_hd__o21ai_1 _08644_ (.A1(_00584_),
    .A2(_02554_),
    .B1(_02558_),
    .Y(_02559_));
 sky130_fd_sc_hd__clkbuf_8 _08645_ (.A(_02525_),
    .X(_02560_));
 sky130_fd_sc_hd__buf_6 _08646_ (.A(_00006_),
    .X(_02561_));
 sky130_fd_sc_hd__buf_6 _08647_ (.A(_02561_),
    .X(_02562_));
 sky130_fd_sc_hd__nand2_1 _08648_ (.A(\H[1][0] ),
    .B(_02562_),
    .Y(_02563_));
 sky130_fd_sc_hd__inv_2 _08649_ (.A(_02563_),
    .Y(_02564_));
 sky130_fd_sc_hd__buf_4 _08650_ (.A(_02562_),
    .X(_02565_));
 sky130_fd_sc_hd__nor2_1 _08651_ (.A(_02565_),
    .B(_02155_),
    .Y(_02566_));
 sky130_fd_sc_hd__buf_6 _08652_ (.A(_02529_),
    .X(_02567_));
 sky130_fd_sc_hd__nand2_1 _08653_ (.A(\H[3][0] ),
    .B(_02567_),
    .Y(_02568_));
 sky130_fd_sc_hd__o211ai_1 _08654_ (.A1(_02567_),
    .A2(_02152_),
    .B1(_02560_),
    .C1(_02568_),
    .Y(_02569_));
 sky130_fd_sc_hd__o31ai_2 _08655_ (.A1(_02560_),
    .A2(_02564_),
    .A3(_02566_),
    .B1(_02569_),
    .Y(_02570_));
 sky130_fd_sc_hd__inv_6 _08656_ (.A(_02555_),
    .Y(_02571_));
 sky130_fd_sc_hd__buf_6 _08657_ (.A(_02571_),
    .X(_02572_));
 sky130_fd_sc_hd__buf_4 _08658_ (.A(_02572_),
    .X(_02573_));
 sky130_fd_sc_hd__a21oi_1 _08659_ (.A1(_02570_),
    .A2(_02573_),
    .B1(_00587_),
    .Y(_02574_));
 sky130_fd_sc_hd__nand2_1 _08660_ (.A(_02559_),
    .B(_02574_),
    .Y(_02575_));
 sky130_fd_sc_hd__nand2_1 _08661_ (.A(\R3[0] ),
    .B(_00587_),
    .Y(_02576_));
 sky130_fd_sc_hd__nand2_2 _08662_ (.A(_02575_),
    .B(_02576_),
    .Y(_02577_));
 sky130_fd_sc_hd__inv_2 _08663_ (.A(_02577_),
    .Y(_02578_));
 sky130_fd_sc_hd__buf_6 _08664_ (.A(_00004_),
    .X(_02579_));
 sky130_fd_sc_hd__inv_4 _08665_ (.A(_02579_),
    .Y(_02580_));
 sky130_fd_sc_hd__buf_6 _08666_ (.A(_02580_),
    .X(_02581_));
 sky130_fd_sc_hd__buf_6 _08667_ (.A(_02581_),
    .X(_02582_));
 sky130_fd_sc_hd__nand2_1 _08668_ (.A(_02582_),
    .B(\Qset[2][0] ),
    .Y(_02583_));
 sky130_fd_sc_hd__buf_4 _08669_ (.A(_00005_),
    .X(_02584_));
 sky130_fd_sc_hd__buf_6 _08670_ (.A(_02579_),
    .X(_02585_));
 sky130_fd_sc_hd__buf_6 _08671_ (.A(_02585_),
    .X(_02586_));
 sky130_fd_sc_hd__nand2_1 _08672_ (.A(_02586_),
    .B(\Qset[3][0] ),
    .Y(_02587_));
 sky130_fd_sc_hd__nand3_1 _08673_ (.A(_02583_),
    .B(_02584_),
    .C(_02587_),
    .Y(_02588_));
 sky130_fd_sc_hd__nand2_1 _08674_ (.A(_02581_),
    .B(\Qset[0][0] ),
    .Y(_02589_));
 sky130_fd_sc_hd__clkinv_4 _08675_ (.A(_00005_),
    .Y(_02590_));
 sky130_fd_sc_hd__buf_4 _08676_ (.A(_02590_),
    .X(_02591_));
 sky130_fd_sc_hd__buf_6 _08677_ (.A(_02579_),
    .X(_02592_));
 sky130_fd_sc_hd__nand2_1 _08678_ (.A(\Qset[1][0] ),
    .B(_02592_),
    .Y(_02593_));
 sky130_fd_sc_hd__nand3_1 _08679_ (.A(_02589_),
    .B(_02591_),
    .C(_02593_),
    .Y(_02594_));
 sky130_fd_sc_hd__nand2_1 _08680_ (.A(_02588_),
    .B(_02594_),
    .Y(_02595_));
 sky130_fd_sc_hd__nand2_1 _08681_ (.A(_02595_),
    .B(_00580_),
    .Y(_02596_));
 sky130_fd_sc_hd__nand2_1 _08682_ (.A(_02138_),
    .B(_02161_),
    .Y(_02597_));
 sky130_fd_sc_hd__nand3_1 _08683_ (.A(_02596_),
    .B(_02597_),
    .C(_02539_),
    .Y(_02598_));
 sky130_fd_sc_hd__nand2_1 _08684_ (.A(_02581_),
    .B(\Oset[2][0] ),
    .Y(_02599_));
 sky130_fd_sc_hd__nand2_1 _08685_ (.A(_02585_),
    .B(\Oset[3][0] ),
    .Y(_02600_));
 sky130_fd_sc_hd__nand3_2 _08686_ (.A(_02599_),
    .B(_00005_),
    .C(_02600_),
    .Y(_02601_));
 sky130_fd_sc_hd__nand2_1 _08687_ (.A(_02581_),
    .B(\Oset[0][0] ),
    .Y(_02602_));
 sky130_fd_sc_hd__nand2_1 _08688_ (.A(_02585_),
    .B(\Oset[1][0] ),
    .Y(_02603_));
 sky130_fd_sc_hd__nand3_4 _08689_ (.A(_02602_),
    .B(_02590_),
    .C(_02603_),
    .Y(_02604_));
 sky130_fd_sc_hd__nand3_1 _08690_ (.A(_02601_),
    .B(_02604_),
    .C(_02551_),
    .Y(_02605_));
 sky130_fd_sc_hd__nand2_1 _08691_ (.A(_02605_),
    .B(_01153_),
    .Y(_02606_));
 sky130_fd_sc_hd__inv_2 _08692_ (.A(_02606_),
    .Y(_02607_));
 sky130_fd_sc_hd__nand2_1 _08693_ (.A(_02598_),
    .B(_02607_),
    .Y(_02608_));
 sky130_fd_sc_hd__a21oi_1 _08694_ (.A1(_02150_),
    .A2(_00583_),
    .B1(_02571_),
    .Y(_02609_));
 sky130_fd_sc_hd__nand2_1 _08695_ (.A(_02608_),
    .B(_02609_),
    .Y(_02610_));
 sky130_fd_sc_hd__buf_6 _08696_ (.A(_02592_),
    .X(_02611_));
 sky130_fd_sc_hd__nor2_1 _08697_ (.A(_02586_),
    .B(_02152_),
    .Y(_02612_));
 sky130_fd_sc_hd__a211o_1 _08698_ (.A1(_02611_),
    .A2(\H[3][0] ),
    .B1(_02591_),
    .C1(_02612_),
    .X(_02613_));
 sky130_fd_sc_hd__nor2_1 _08699_ (.A(_02586_),
    .B(_02155_),
    .Y(_02614_));
 sky130_fd_sc_hd__a211o_1 _08700_ (.A1(_02586_),
    .A2(\H[1][0] ),
    .B1(_02584_),
    .C1(_02614_),
    .X(_02615_));
 sky130_fd_sc_hd__nand3_1 _08701_ (.A(_02613_),
    .B(_02615_),
    .C(_02571_),
    .Y(_02616_));
 sky130_fd_sc_hd__nand2_1 _08702_ (.A(_02610_),
    .B(_02616_),
    .Y(_02617_));
 sky130_fd_sc_hd__nand2_1 _08703_ (.A(_02617_),
    .B(_01551_),
    .Y(_02618_));
 sky130_fd_sc_hd__nand2_4 _08704_ (.A(_02618_),
    .B(_02158_),
    .Y(_02619_));
 sky130_fd_sc_hd__buf_6 _08705_ (.A(_02619_),
    .X(_02620_));
 sky130_fd_sc_hd__nand2_2 _08706_ (.A(_02620_),
    .B(_02577_),
    .Y(_02621_));
 sky130_fd_sc_hd__o21ai_4 _08707_ (.A1(_00622_),
    .A2(_02578_),
    .B1(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__xor2_4 _08708_ (.A(_02160_),
    .B(_02622_),
    .X(_02623_));
 sky130_fd_sc_hd__clkbuf_4 _08709_ (.A(_00000_),
    .X(_02624_));
 sky130_fd_sc_hd__clkbuf_4 _08710_ (.A(_02624_),
    .X(_02625_));
 sky130_fd_sc_hd__inv_2 _08711_ (.A(_00001_),
    .Y(_02626_));
 sky130_fd_sc_hd__nor2_1 _08712_ (.A(_02625_),
    .B(_02152_),
    .Y(_02627_));
 sky130_fd_sc_hd__a211o_1 _08713_ (.A1(\H[3][0] ),
    .A2(_02625_),
    .B1(_02626_),
    .C1(_02627_),
    .X(_02628_));
 sky130_fd_sc_hd__nor2_1 _08714_ (.A(_02625_),
    .B(_02155_),
    .Y(_02629_));
 sky130_fd_sc_hd__a211o_1 _08715_ (.A1(\H[1][0] ),
    .A2(_02625_),
    .B1(_00001_),
    .C1(_02629_),
    .X(_02630_));
 sky130_fd_sc_hd__mux2_1 _08716_ (.A0(\Qset[2][0] ),
    .A1(\Qset[3][0] ),
    .S(_00000_),
    .X(_02631_));
 sky130_fd_sc_hd__inv_2 _08717_ (.A(_02624_),
    .Y(_02632_));
 sky130_fd_sc_hd__a21o_1 _08718_ (.A1(\Qset[1][0] ),
    .A2(_02624_),
    .B1(_00001_),
    .X(_02633_));
 sky130_fd_sc_hd__a21o_1 _08719_ (.A1(\Qset[0][0] ),
    .A2(_02632_),
    .B1(_02633_),
    .X(_02634_));
 sky130_fd_sc_hd__o21a_1 _08720_ (.A1(_02626_),
    .A2(_02631_),
    .B1(_02634_),
    .X(_02635_));
 sky130_fd_sc_hd__nor2_1 _08721_ (.A(_02624_),
    .B(_02142_),
    .Y(_02636_));
 sky130_fd_sc_hd__a211o_1 _08722_ (.A1(\Oset[3][0] ),
    .A2(_02624_),
    .B1(_02626_),
    .C1(_02636_),
    .X(_02637_));
 sky130_fd_sc_hd__nor2_1 _08723_ (.A(_02624_),
    .B(_02146_),
    .Y(_02638_));
 sky130_fd_sc_hd__a211o_1 _08724_ (.A1(\Oset[1][0] ),
    .A2(_02624_),
    .B1(_00001_),
    .C1(_02638_),
    .X(_02639_));
 sky130_fd_sc_hd__a21o_1 _08725_ (.A1(_02637_),
    .A2(_02639_),
    .B1(_00646_),
    .X(_02640_));
 sky130_fd_sc_hd__o211a_1 _08726_ (.A1(Oreg3),
    .A2(_02635_),
    .B1(_00626_),
    .C1(_02640_),
    .X(_02641_));
 sky130_fd_sc_hd__a311o_1 _08727_ (.A1(_01536_),
    .A2(_02628_),
    .A3(_02630_),
    .B1(_00548_),
    .C1(_02641_),
    .X(_02642_));
 sky130_fd_sc_hd__o21ai_2 _08728_ (.A1(_00622_),
    .A2(_02620_),
    .B1(_02642_),
    .Y(_02643_));
 sky130_fd_sc_hd__xor2_2 _08729_ (.A(_00832_),
    .B(_02643_),
    .X(_02644_));
 sky130_fd_sc_hd__xor2_4 _08730_ (.A(_02623_),
    .B(_02644_),
    .X(_02645_));
 sky130_fd_sc_hd__inv_2 _08731_ (.A(_02645_),
    .Y(_02646_));
 sky130_fd_sc_hd__nand2_1 _08732_ (.A(CMD_addition),
    .B(\current_state[6] ),
    .Y(_02647_));
 sky130_fd_sc_hd__inv_2 _08733_ (.A(_02647_),
    .Y(_02648_));
 sky130_fd_sc_hd__buf_4 _08734_ (.A(_02648_),
    .X(_02649_));
 sky130_fd_sc_hd__buf_6 _08735_ (.A(_00635_),
    .X(_02650_));
 sky130_fd_sc_hd__nor2_1 _08736_ (.A(\result_reg_add[0] ),
    .B(_02648_),
    .Y(_02651_));
 sky130_fd_sc_hd__a211o_1 _08737_ (.A1(_02646_),
    .A2(_02649_),
    .B1(_02650_),
    .C1(_02651_),
    .X(_02652_));
 sky130_fd_sc_hd__inv_2 _08738_ (.A(_02652_),
    .Y(_00244_));
 sky130_fd_sc_hd__clkbuf_4 _08739_ (.A(_02647_),
    .X(_02653_));
 sky130_fd_sc_hd__clkbuf_4 _08740_ (.A(_02653_),
    .X(_02654_));
 sky130_fd_sc_hd__nand2_1 _08741_ (.A(_02581_),
    .B(\Qset[2][1] ),
    .Y(_02655_));
 sky130_fd_sc_hd__nand2_1 _08742_ (.A(_02585_),
    .B(\Qset[3][1] ),
    .Y(_02656_));
 sky130_fd_sc_hd__nand3_1 _08743_ (.A(_02655_),
    .B(_00005_),
    .C(_02656_),
    .Y(_02657_));
 sky130_fd_sc_hd__nand2_1 _08744_ (.A(_02581_),
    .B(\Qset[0][1] ),
    .Y(_02658_));
 sky130_fd_sc_hd__nand2_1 _08745_ (.A(_02585_),
    .B(\Qset[1][1] ),
    .Y(_02659_));
 sky130_fd_sc_hd__nand3_1 _08746_ (.A(_02658_),
    .B(_02590_),
    .C(_02659_),
    .Y(_02660_));
 sky130_fd_sc_hd__nand2_2 _08747_ (.A(_02657_),
    .B(_02660_),
    .Y(_02661_));
 sky130_fd_sc_hd__nand2_1 _08748_ (.A(_02661_),
    .B(_00580_),
    .Y(_02662_));
 sky130_fd_sc_hd__nand2_1 _08749_ (.A(_02178_),
    .B(\shift.Q ),
    .Y(_02663_));
 sky130_fd_sc_hd__nand3_1 _08750_ (.A(_02662_),
    .B(_02663_),
    .C(_02539_),
    .Y(_02664_));
 sky130_fd_sc_hd__nand2_1 _08751_ (.A(_02580_),
    .B(\Oset[2][1] ),
    .Y(_02665_));
 sky130_fd_sc_hd__nand2_1 _08752_ (.A(_02579_),
    .B(\Oset[3][1] ),
    .Y(_02666_));
 sky130_fd_sc_hd__nand3_2 _08753_ (.A(_02665_),
    .B(_00005_),
    .C(_02666_),
    .Y(_02667_));
 sky130_fd_sc_hd__nand2_1 _08754_ (.A(_02580_),
    .B(\Oset[0][1] ),
    .Y(_02668_));
 sky130_fd_sc_hd__nand2_1 _08755_ (.A(_02579_),
    .B(\Oset[1][1] ),
    .Y(_02669_));
 sky130_fd_sc_hd__nand3_2 _08756_ (.A(_02668_),
    .B(_02590_),
    .C(_02669_),
    .Y(_02670_));
 sky130_fd_sc_hd__nand3_1 _08757_ (.A(_02667_),
    .B(_02670_),
    .C(_02551_),
    .Y(_02671_));
 sky130_fd_sc_hd__nand2_1 _08758_ (.A(_02671_),
    .B(_01153_),
    .Y(_02672_));
 sky130_fd_sc_hd__inv_2 _08759_ (.A(_02672_),
    .Y(_02673_));
 sky130_fd_sc_hd__nand2_1 _08760_ (.A(_02664_),
    .B(_02673_),
    .Y(_02674_));
 sky130_fd_sc_hd__a21oi_1 _08761_ (.A1(_02185_),
    .A2(_00583_),
    .B1(_02571_),
    .Y(_02675_));
 sky130_fd_sc_hd__nand2_1 _08762_ (.A(_02674_),
    .B(_02675_),
    .Y(_02676_));
 sky130_fd_sc_hd__nor2_1 _08763_ (.A(_02579_),
    .B(_02189_),
    .Y(_02677_));
 sky130_fd_sc_hd__a211o_1 _08764_ (.A1(_02585_),
    .A2(\H[1][1] ),
    .B1(_00005_),
    .C1(_02677_),
    .X(_02678_));
 sky130_fd_sc_hd__nor2_1 _08765_ (.A(_02579_),
    .B(_02186_),
    .Y(_02679_));
 sky130_fd_sc_hd__a211o_1 _08766_ (.A1(_02585_),
    .A2(\H[3][1] ),
    .B1(_02590_),
    .C1(_02679_),
    .X(_02680_));
 sky130_fd_sc_hd__nand2_1 _08767_ (.A(_02678_),
    .B(_02680_),
    .Y(_02681_));
 sky130_fd_sc_hd__inv_2 _08768_ (.A(_02681_),
    .Y(_02682_));
 sky130_fd_sc_hd__nand2_1 _08769_ (.A(_02682_),
    .B(_02571_),
    .Y(_02683_));
 sky130_fd_sc_hd__nand2_1 _08770_ (.A(_02676_),
    .B(_02683_),
    .Y(_02684_));
 sky130_fd_sc_hd__nand2_1 _08771_ (.A(_02684_),
    .B(_01551_),
    .Y(_02685_));
 sky130_fd_sc_hd__nand2_1 _08772_ (.A(_02685_),
    .B(_02192_),
    .Y(_02686_));
 sky130_fd_sc_hd__buf_4 _08773_ (.A(_02686_),
    .X(_02687_));
 sky130_fd_sc_hd__clkbuf_4 _08774_ (.A(_02625_),
    .X(_02688_));
 sky130_fd_sc_hd__nor2_1 _08775_ (.A(_02688_),
    .B(_02186_),
    .Y(_02689_));
 sky130_fd_sc_hd__a211o_1 _08776_ (.A1(\H[3][1] ),
    .A2(_02688_),
    .B1(_02626_),
    .C1(_02689_),
    .X(_02690_));
 sky130_fd_sc_hd__nor2_1 _08777_ (.A(_02688_),
    .B(_02189_),
    .Y(_02691_));
 sky130_fd_sc_hd__a211o_1 _08778_ (.A1(\H[1][1] ),
    .A2(_02688_),
    .B1(_00001_),
    .C1(_02691_),
    .X(_02692_));
 sky130_fd_sc_hd__mux2_1 _08779_ (.A0(\Qset[2][1] ),
    .A1(\Qset[3][1] ),
    .S(_02624_),
    .X(_02693_));
 sky130_fd_sc_hd__a21o_1 _08780_ (.A1(\Qset[1][1] ),
    .A2(_02624_),
    .B1(_00001_),
    .X(_02694_));
 sky130_fd_sc_hd__a21o_1 _08781_ (.A1(\Qset[0][1] ),
    .A2(_02632_),
    .B1(_02694_),
    .X(_02695_));
 sky130_fd_sc_hd__o21a_1 _08782_ (.A1(_02626_),
    .A2(_02693_),
    .B1(_02695_),
    .X(_02696_));
 sky130_fd_sc_hd__nor2_1 _08783_ (.A(_02625_),
    .B(_02179_),
    .Y(_02697_));
 sky130_fd_sc_hd__a211o_1 _08784_ (.A1(\Oset[3][1] ),
    .A2(_02625_),
    .B1(_02626_),
    .C1(_02697_),
    .X(_02698_));
 sky130_fd_sc_hd__nor2_1 _08785_ (.A(_02624_),
    .B(_02182_),
    .Y(_02699_));
 sky130_fd_sc_hd__a211o_1 _08786_ (.A1(\Oset[1][1] ),
    .A2(_02625_),
    .B1(_00001_),
    .C1(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__a21o_1 _08787_ (.A1(_02698_),
    .A2(_02700_),
    .B1(_00646_),
    .X(_02701_));
 sky130_fd_sc_hd__o211a_1 _08788_ (.A1(Oreg3),
    .A2(_02696_),
    .B1(_00626_),
    .C1(_02701_),
    .X(_02702_));
 sky130_fd_sc_hd__a311o_1 _08789_ (.A1(_01536_),
    .A2(_02690_),
    .A3(_02692_),
    .B1(_00548_),
    .C1(_02702_),
    .X(_02703_));
 sky130_fd_sc_hd__o21ai_1 _08790_ (.A1(_00622_),
    .A2(_02687_),
    .B1(_02703_),
    .Y(_02704_));
 sky130_fd_sc_hd__nand2_1 _08791_ (.A(_02522_),
    .B(\Qset[2][1] ),
    .Y(_02705_));
 sky130_fd_sc_hd__nand2_1 _08792_ (.A(_02527_),
    .B(\Qset[3][1] ),
    .Y(_02706_));
 sky130_fd_sc_hd__nand3_1 _08793_ (.A(_02705_),
    .B(_00007_),
    .C(_02706_),
    .Y(_02707_));
 sky130_fd_sc_hd__nand2_1 _08794_ (.A(_02522_),
    .B(\Qset[0][1] ),
    .Y(_02708_));
 sky130_fd_sc_hd__nand2_1 _08795_ (.A(_02527_),
    .B(\Qset[1][1] ),
    .Y(_02709_));
 sky130_fd_sc_hd__nand3_1 _08796_ (.A(_02708_),
    .B(_02533_),
    .C(_02709_),
    .Y(_02710_));
 sky130_fd_sc_hd__nand2_2 _08797_ (.A(_02707_),
    .B(_02710_),
    .Y(_02711_));
 sky130_fd_sc_hd__o21ai_1 _08798_ (.A1(_00580_),
    .A2(_00669_),
    .B1(_02539_),
    .Y(_02712_));
 sky130_fd_sc_hd__inv_2 _08799_ (.A(_02712_),
    .Y(_02713_));
 sky130_fd_sc_hd__o21ai_1 _08800_ (.A1(_02161_),
    .A2(_02711_),
    .B1(_02713_),
    .Y(_02714_));
 sky130_fd_sc_hd__nand2_1 _08801_ (.A(_02527_),
    .B(\Oset[1][1] ),
    .Y(_02715_));
 sky130_fd_sc_hd__o211ai_1 _08802_ (.A1(_02527_),
    .A2(_02182_),
    .B1(_02534_),
    .C1(_02715_),
    .Y(_02716_));
 sky130_fd_sc_hd__nand2_1 _08803_ (.A(_02527_),
    .B(\Oset[3][1] ),
    .Y(_02717_));
 sky130_fd_sc_hd__o211ai_1 _08804_ (.A1(_02527_),
    .A2(_02179_),
    .B1(_00007_),
    .C1(_02717_),
    .Y(_02718_));
 sky130_fd_sc_hd__nand2_2 _08805_ (.A(_02716_),
    .B(_02718_),
    .Y(_02719_));
 sky130_fd_sc_hd__nand2_1 _08806_ (.A(_02719_),
    .B(_02551_),
    .Y(_02720_));
 sky130_fd_sc_hd__nand3_1 _08807_ (.A(_02714_),
    .B(_02720_),
    .C(_01154_),
    .Y(_02721_));
 sky130_fd_sc_hd__o21ai_1 _08808_ (.A1(_01153_),
    .A2(_00669_),
    .B1(_02555_),
    .Y(_02722_));
 sky130_fd_sc_hd__inv_2 _08809_ (.A(_02722_),
    .Y(_02723_));
 sky130_fd_sc_hd__nand2_1 _08810_ (.A(_02721_),
    .B(_02723_),
    .Y(_02724_));
 sky130_fd_sc_hd__nand2_1 _08811_ (.A(_02527_),
    .B(\H[3][1] ),
    .Y(_02725_));
 sky130_fd_sc_hd__o21ai_1 _08812_ (.A1(_02561_),
    .A2(_02186_),
    .B1(_02725_),
    .Y(_02726_));
 sky130_fd_sc_hd__buf_4 _08813_ (.A(_00007_),
    .X(_02727_));
 sky130_fd_sc_hd__o21a_1 _08814_ (.A1(\H[1][1] ),
    .A2(_02522_),
    .B1(_02534_),
    .X(_02728_));
 sky130_fd_sc_hd__nand2_1 _08815_ (.A(_02522_),
    .B(_02189_),
    .Y(_02729_));
 sky130_fd_sc_hd__a22oi_4 _08816_ (.A1(_02726_),
    .A2(_02727_),
    .B1(_02728_),
    .B2(_02729_),
    .Y(_02730_));
 sky130_fd_sc_hd__a21oi_1 _08817_ (.A1(_02730_),
    .A2(_02571_),
    .B1(_00586_),
    .Y(_02731_));
 sky130_fd_sc_hd__nand2_1 _08818_ (.A(_02724_),
    .B(_02731_),
    .Y(_02732_));
 sky130_fd_sc_hd__nand2_1 _08819_ (.A(_00586_),
    .B(\R3[1] ),
    .Y(_02733_));
 sky130_fd_sc_hd__nand2_2 _08820_ (.A(_02732_),
    .B(_02733_),
    .Y(_02734_));
 sky130_fd_sc_hd__inv_2 _08821_ (.A(_02734_),
    .Y(_02735_));
 sky130_fd_sc_hd__nand2_1 _08822_ (.A(_02687_),
    .B(_02734_),
    .Y(_02736_));
 sky130_fd_sc_hd__or2_1 _08823_ (.A(_02736_),
    .B(_02621_),
    .X(_02737_));
 sky130_fd_sc_hd__inv_2 _08824_ (.A(_02686_),
    .Y(_02738_));
 sky130_fd_sc_hd__nand2_1 _08825_ (.A(_02620_),
    .B(_02734_),
    .Y(_02739_));
 sky130_fd_sc_hd__o21ai_1 _08826_ (.A1(_02578_),
    .A2(_02738_),
    .B1(_02739_),
    .Y(_02740_));
 sky130_fd_sc_hd__nand3_1 _08827_ (.A(_02737_),
    .B(_00622_),
    .C(_02740_),
    .Y(_02741_));
 sky130_fd_sc_hd__o21ai_1 _08828_ (.A1(_00622_),
    .A2(_02735_),
    .B1(_02741_),
    .Y(_02742_));
 sky130_fd_sc_hd__xor2_1 _08829_ (.A(_00536_),
    .B(_02742_),
    .X(_02743_));
 sky130_fd_sc_hd__or2_1 _08830_ (.A(_02704_),
    .B(_02743_),
    .X(_02744_));
 sky130_fd_sc_hd__nand2_1 _08831_ (.A(_02743_),
    .B(_02704_),
    .Y(_02745_));
 sky130_fd_sc_hd__mux2_1 _08832_ (.A0(_00536_),
    .A1(_02643_),
    .S(_02622_),
    .X(_02746_));
 sky130_fd_sc_hd__inv_2 _08833_ (.A(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__a21o_1 _08834_ (.A1(_02744_),
    .A2(_02745_),
    .B1(_02747_),
    .X(_02748_));
 sky130_fd_sc_hd__nand3_1 _08835_ (.A(_02747_),
    .B(_02744_),
    .C(_02745_),
    .Y(_02749_));
 sky130_fd_sc_hd__and2_2 _08836_ (.A(_02748_),
    .B(_02749_),
    .X(_02750_));
 sky130_fd_sc_hd__nor2_1 _08837_ (.A(_02653_),
    .B(_02750_),
    .Y(_02751_));
 sky130_fd_sc_hd__a211o_1 _08838_ (.A1(_00703_),
    .A2(_02654_),
    .B1(_02650_),
    .C1(_02751_),
    .X(_02752_));
 sky130_fd_sc_hd__inv_2 _08839_ (.A(_02752_),
    .Y(_00245_));
 sky130_fd_sc_hd__clkbuf_4 _08840_ (.A(_00635_),
    .X(_02753_));
 sky130_fd_sc_hd__nand2_1 _08841_ (.A(_02581_),
    .B(\Qset[2][2] ),
    .Y(_02754_));
 sky130_fd_sc_hd__nand2_1 _08842_ (.A(_02592_),
    .B(\Qset[3][2] ),
    .Y(_02755_));
 sky130_fd_sc_hd__nand3_1 _08843_ (.A(_02754_),
    .B(_02584_),
    .C(_02755_),
    .Y(_02756_));
 sky130_fd_sc_hd__nand2_1 _08844_ (.A(_02581_),
    .B(\Qset[0][2] ),
    .Y(_02757_));
 sky130_fd_sc_hd__nand2_1 _08845_ (.A(_02585_),
    .B(\Qset[1][2] ),
    .Y(_02758_));
 sky130_fd_sc_hd__nand3_1 _08846_ (.A(_02757_),
    .B(_02590_),
    .C(_02758_),
    .Y(_02759_));
 sky130_fd_sc_hd__nand2_2 _08847_ (.A(_02756_),
    .B(_02759_),
    .Y(_02760_));
 sky130_fd_sc_hd__nand2_1 _08848_ (.A(_02760_),
    .B(_00580_),
    .Y(_02761_));
 sky130_fd_sc_hd__nand2_1 _08849_ (.A(_02201_),
    .B(_02161_),
    .Y(_02762_));
 sky130_fd_sc_hd__nand3_1 _08850_ (.A(_02761_),
    .B(_02762_),
    .C(_02539_),
    .Y(_02763_));
 sky130_fd_sc_hd__nand2_1 _08851_ (.A(_02580_),
    .B(\Oset[2][2] ),
    .Y(_02764_));
 sky130_fd_sc_hd__nand2_1 _08852_ (.A(_02585_),
    .B(\Oset[3][2] ),
    .Y(_02765_));
 sky130_fd_sc_hd__nand3_1 _08853_ (.A(_02764_),
    .B(_00005_),
    .C(_02765_),
    .Y(_02766_));
 sky130_fd_sc_hd__nand2_1 _08854_ (.A(_02580_),
    .B(\Oset[0][2] ),
    .Y(_02767_));
 sky130_fd_sc_hd__nand2_1 _08855_ (.A(_02579_),
    .B(\Oset[1][2] ),
    .Y(_02768_));
 sky130_fd_sc_hd__nand3_2 _08856_ (.A(_02767_),
    .B(_02590_),
    .C(_02768_),
    .Y(_02769_));
 sky130_fd_sc_hd__nand3_1 _08857_ (.A(_02766_),
    .B(_02769_),
    .C(_02551_),
    .Y(_02770_));
 sky130_fd_sc_hd__nand2_1 _08858_ (.A(_02770_),
    .B(_01153_),
    .Y(_02771_));
 sky130_fd_sc_hd__inv_2 _08859_ (.A(_02771_),
    .Y(_02772_));
 sky130_fd_sc_hd__nand2_1 _08860_ (.A(_02763_),
    .B(_02772_),
    .Y(_02773_));
 sky130_fd_sc_hd__nand2_1 _08861_ (.A(_02206_),
    .B(_00583_),
    .Y(_02774_));
 sky130_fd_sc_hd__nand2_1 _08862_ (.A(_02773_),
    .B(_02774_),
    .Y(_02775_));
 sky130_fd_sc_hd__nand2_1 _08863_ (.A(_02775_),
    .B(_02555_),
    .Y(_02776_));
 sky130_fd_sc_hd__nor2_1 _08864_ (.A(_02592_),
    .B(_02207_),
    .Y(_02777_));
 sky130_fd_sc_hd__a211o_1 _08865_ (.A1(_02586_),
    .A2(\H[3][2] ),
    .B1(_02591_),
    .C1(_02777_),
    .X(_02778_));
 sky130_fd_sc_hd__nor2_1 _08866_ (.A(_02592_),
    .B(_02210_),
    .Y(_02779_));
 sky130_fd_sc_hd__a211o_1 _08867_ (.A1(_02586_),
    .A2(\H[1][2] ),
    .B1(_02584_),
    .C1(_02779_),
    .X(_02780_));
 sky130_fd_sc_hd__nand2_2 _08868_ (.A(_02778_),
    .B(_02780_),
    .Y(_02781_));
 sky130_fd_sc_hd__a21oi_1 _08869_ (.A1(_02781_),
    .A2(_02571_),
    .B1(_00586_),
    .Y(_02782_));
 sky130_fd_sc_hd__nand2_1 _08870_ (.A(_02776_),
    .B(_02782_),
    .Y(_02783_));
 sky130_fd_sc_hd__nand2_2 _08871_ (.A(_02783_),
    .B(_02213_),
    .Y(_02784_));
 sky130_fd_sc_hd__buf_6 _08872_ (.A(_02784_),
    .X(_02785_));
 sky130_fd_sc_hd__and2_1 _08873_ (.A(_02785_),
    .B(_02577_),
    .X(_02786_));
 sky130_fd_sc_hd__buf_6 _08874_ (.A(_02522_),
    .X(_02787_));
 sky130_fd_sc_hd__nand2_1 _08875_ (.A(_02787_),
    .B(\Qset[2][2] ),
    .Y(_02788_));
 sky130_fd_sc_hd__nand2_1 _08876_ (.A(_02562_),
    .B(\Qset[3][2] ),
    .Y(_02789_));
 sky130_fd_sc_hd__nand3_2 _08877_ (.A(_02788_),
    .B(_02525_),
    .C(_02789_),
    .Y(_02790_));
 sky130_fd_sc_hd__nand2_1 _08878_ (.A(_02787_),
    .B(\Qset[0][2] ),
    .Y(_02791_));
 sky130_fd_sc_hd__nand2_1 _08879_ (.A(_02562_),
    .B(\Qset[1][2] ),
    .Y(_02792_));
 sky130_fd_sc_hd__nand3_2 _08880_ (.A(_02791_),
    .B(_02535_),
    .C(_02792_),
    .Y(_02793_));
 sky130_fd_sc_hd__nand3_1 _08881_ (.A(_02790_),
    .B(_02793_),
    .C(_00581_),
    .Y(_02794_));
 sky130_fd_sc_hd__o21ai_1 _08882_ (.A1(_00681_),
    .A2(_00580_),
    .B1(_02539_),
    .Y(_02795_));
 sky130_fd_sc_hd__inv_2 _08883_ (.A(_02795_),
    .Y(_02796_));
 sky130_fd_sc_hd__nand2_1 _08884_ (.A(_02794_),
    .B(_02796_),
    .Y(_02797_));
 sky130_fd_sc_hd__buf_6 _08885_ (.A(_02561_),
    .X(_02798_));
 sky130_fd_sc_hd__nand2_1 _08886_ (.A(_02798_),
    .B(\Oset[1][2] ),
    .Y(_02799_));
 sky130_fd_sc_hd__buf_6 _08887_ (.A(_02534_),
    .X(_02800_));
 sky130_fd_sc_hd__nand2_1 _08888_ (.A(_02799_),
    .B(_02800_),
    .Y(_02801_));
 sky130_fd_sc_hd__nand2_1 _08889_ (.A(_02522_),
    .B(\Oset[0][2] ),
    .Y(_02802_));
 sky130_fd_sc_hd__inv_2 _08890_ (.A(_02802_),
    .Y(_02803_));
 sky130_fd_sc_hd__nand2_1 _08891_ (.A(_02787_),
    .B(\Oset[2][2] ),
    .Y(_02804_));
 sky130_fd_sc_hd__nand2_1 _08892_ (.A(_02798_),
    .B(\Oset[3][2] ),
    .Y(_02805_));
 sky130_fd_sc_hd__nand3_1 _08893_ (.A(_02804_),
    .B(_02525_),
    .C(_02805_),
    .Y(_02806_));
 sky130_fd_sc_hd__o21ai_4 _08894_ (.A1(_02801_),
    .A2(_02803_),
    .B1(_02806_),
    .Y(_02807_));
 sky130_fd_sc_hd__nand2_1 _08895_ (.A(_02807_),
    .B(_02552_),
    .Y(_02808_));
 sky130_fd_sc_hd__nand3_1 _08896_ (.A(_02797_),
    .B(_02808_),
    .C(_01155_),
    .Y(_02809_));
 sky130_fd_sc_hd__o21ai_1 _08897_ (.A1(_00681_),
    .A2(_01154_),
    .B1(_02555_),
    .Y(_02810_));
 sky130_fd_sc_hd__inv_2 _08898_ (.A(_02810_),
    .Y(_02811_));
 sky130_fd_sc_hd__nand2_1 _08899_ (.A(_02809_),
    .B(_02811_),
    .Y(_02812_));
 sky130_fd_sc_hd__nor2_1 _08900_ (.A(_02529_),
    .B(_02210_),
    .Y(_02813_));
 sky130_fd_sc_hd__a21o_1 _08901_ (.A1(_02798_),
    .A2(\H[1][2] ),
    .B1(_02525_),
    .X(_02814_));
 sky130_fd_sc_hd__nand2_1 _08902_ (.A(_02545_),
    .B(\H[3][2] ),
    .Y(_02815_));
 sky130_fd_sc_hd__o211ai_1 _08903_ (.A1(_02529_),
    .A2(_02207_),
    .B1(_02526_),
    .C1(_02815_),
    .Y(_02816_));
 sky130_fd_sc_hd__o21ai_2 _08904_ (.A1(_02813_),
    .A2(_02814_),
    .B1(_02816_),
    .Y(_02817_));
 sky130_fd_sc_hd__a21oi_1 _08905_ (.A1(_02817_),
    .A2(_02572_),
    .B1(_00586_),
    .Y(_02818_));
 sky130_fd_sc_hd__nand2_1 _08906_ (.A(_02812_),
    .B(_02818_),
    .Y(_02819_));
 sky130_fd_sc_hd__nand2_1 _08907_ (.A(\R2[0] ),
    .B(_00587_),
    .Y(_02820_));
 sky130_fd_sc_hd__nand2_4 _08908_ (.A(_02819_),
    .B(_02820_),
    .Y(_02821_));
 sky130_fd_sc_hd__nand2_1 _08909_ (.A(_02687_),
    .B(_02821_),
    .Y(_02822_));
 sky130_fd_sc_hd__nand2_1 _08910_ (.A(_02619_),
    .B(_02821_),
    .Y(_02823_));
 sky130_fd_sc_hd__nand2_1 _08911_ (.A(_02736_),
    .B(_02823_),
    .Y(_02824_));
 sky130_fd_sc_hd__o21a_1 _08912_ (.A1(_02739_),
    .A2(_02822_),
    .B1(_02824_),
    .X(_02825_));
 sky130_fd_sc_hd__or2_1 _08913_ (.A(_02786_),
    .B(_02825_),
    .X(_02826_));
 sky130_fd_sc_hd__nand2_1 _08914_ (.A(_02825_),
    .B(_02786_),
    .Y(_02827_));
 sky130_fd_sc_hd__nand3b_2 _08915_ (.A_N(_02737_),
    .B(_02826_),
    .C(_02827_),
    .Y(_02828_));
 sky130_fd_sc_hd__xnor2_1 _08916_ (.A(_02786_),
    .B(_02825_),
    .Y(_02829_));
 sky130_fd_sc_hd__nand2_1 _08917_ (.A(_02829_),
    .B(_02737_),
    .Y(_02830_));
 sky130_fd_sc_hd__nand3_1 _08918_ (.A(_02828_),
    .B(_02830_),
    .C(_00622_),
    .Y(_02831_));
 sky130_fd_sc_hd__nand2_1 _08919_ (.A(_02821_),
    .B(_00549_),
    .Y(_02832_));
 sky130_fd_sc_hd__a21o_1 _08920_ (.A1(_02831_),
    .A2(_02832_),
    .B1(_00536_),
    .X(_02833_));
 sky130_fd_sc_hd__nand3_1 _08921_ (.A(_02831_),
    .B(_00536_),
    .C(_02832_),
    .Y(_02834_));
 sky130_fd_sc_hd__nand2_1 _08922_ (.A(_02833_),
    .B(_02834_),
    .Y(_02835_));
 sky130_fd_sc_hd__clkbuf_4 _08923_ (.A(_02688_),
    .X(_02836_));
 sky130_fd_sc_hd__clkbuf_4 _08924_ (.A(_02626_),
    .X(_02837_));
 sky130_fd_sc_hd__nor2_1 _08925_ (.A(_02688_),
    .B(_02207_),
    .Y(_02838_));
 sky130_fd_sc_hd__a211o_1 _08926_ (.A1(\H[3][2] ),
    .A2(_02836_),
    .B1(_02837_),
    .C1(_02838_),
    .X(_02839_));
 sky130_fd_sc_hd__buf_4 _08927_ (.A(_00001_),
    .X(_02840_));
 sky130_fd_sc_hd__nor2_1 _08928_ (.A(_02688_),
    .B(_02210_),
    .Y(_02841_));
 sky130_fd_sc_hd__a211o_1 _08929_ (.A1(\H[1][2] ),
    .A2(_02836_),
    .B1(_02840_),
    .C1(_02841_),
    .X(_02842_));
 sky130_fd_sc_hd__mux2_1 _08930_ (.A0(\Oset[2][2] ),
    .A1(\Oset[3][2] ),
    .S(_02688_),
    .X(_02843_));
 sky130_fd_sc_hd__a21o_1 _08931_ (.A1(\Oset[1][2] ),
    .A2(_02688_),
    .B1(_02840_),
    .X(_02844_));
 sky130_fd_sc_hd__a21o_1 _08932_ (.A1(\Oset[0][2] ),
    .A2(_02632_),
    .B1(_02844_),
    .X(_02845_));
 sky130_fd_sc_hd__o21ai_1 _08933_ (.A1(_02837_),
    .A2(_02843_),
    .B1(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hd__mux2_1 _08934_ (.A0(\Qset[2][2] ),
    .A1(\Qset[3][2] ),
    .S(_02625_),
    .X(_02847_));
 sky130_fd_sc_hd__a21o_1 _08935_ (.A1(\Qset[1][2] ),
    .A2(_02625_),
    .B1(_00001_),
    .X(_02848_));
 sky130_fd_sc_hd__a21o_1 _08936_ (.A1(\Qset[0][2] ),
    .A2(_02632_),
    .B1(_02848_),
    .X(_02849_));
 sky130_fd_sc_hd__o21ai_1 _08937_ (.A1(_02837_),
    .A2(_02847_),
    .B1(_02849_),
    .Y(_02850_));
 sky130_fd_sc_hd__a21o_1 _08938_ (.A1(_02850_),
    .A2(_00646_),
    .B1(_01536_),
    .X(_02851_));
 sky130_fd_sc_hd__a21oi_1 _08939_ (.A1(_00621_),
    .A2(_02846_),
    .B1(_02851_),
    .Y(_02852_));
 sky130_fd_sc_hd__a311o_1 _08940_ (.A1(_01536_),
    .A2(_02839_),
    .A3(_02842_),
    .B1(_00548_),
    .C1(_02852_),
    .X(_02853_));
 sky130_fd_sc_hd__o21ai_1 _08941_ (.A1(_00622_),
    .A2(_02785_),
    .B1(_02853_),
    .Y(_02854_));
 sky130_fd_sc_hd__nand2_1 _08942_ (.A(_02835_),
    .B(_02854_),
    .Y(_02855_));
 sky130_fd_sc_hd__nand3b_1 _08943_ (.A_N(_02854_),
    .B(_02833_),
    .C(_02834_),
    .Y(_02856_));
 sky130_fd_sc_hd__nand2_1 _08944_ (.A(_02749_),
    .B(_02744_),
    .Y(_02857_));
 sky130_fd_sc_hd__a21o_1 _08945_ (.A1(_02855_),
    .A2(_02856_),
    .B1(_02857_),
    .X(_02858_));
 sky130_fd_sc_hd__nand3_1 _08946_ (.A(_02857_),
    .B(_02855_),
    .C(_02856_),
    .Y(_02859_));
 sky130_fd_sc_hd__and2_2 _08947_ (.A(_02858_),
    .B(_02859_),
    .X(_02860_));
 sky130_fd_sc_hd__nor2_1 _08948_ (.A(_02653_),
    .B(_02860_),
    .Y(_02861_));
 sky130_fd_sc_hd__a211o_1 _08949_ (.A1(_00729_),
    .A2(_02654_),
    .B1(_02753_),
    .C1(_02861_),
    .X(_02862_));
 sky130_fd_sc_hd__inv_2 _08950_ (.A(_02862_),
    .Y(_00246_));
 sky130_fd_sc_hd__nor2_1 _08951_ (.A(_02737_),
    .B(_02829_),
    .Y(_02863_));
 sky130_fd_sc_hd__nand2_1 _08952_ (.A(_02787_),
    .B(\Qset[2][3] ),
    .Y(_02864_));
 sky130_fd_sc_hd__nand2_1 _08953_ (.A(_02544_),
    .B(\Qset[3][3] ),
    .Y(_02865_));
 sky130_fd_sc_hd__nand3_1 _08954_ (.A(_02864_),
    .B(_02525_),
    .C(_02865_),
    .Y(_02866_));
 sky130_fd_sc_hd__nand2_1 _08955_ (.A(_02522_),
    .B(\Qset[0][3] ),
    .Y(_02867_));
 sky130_fd_sc_hd__nand2_1 _08956_ (.A(_02528_),
    .B(\Qset[1][3] ),
    .Y(_02868_));
 sky130_fd_sc_hd__nand3_1 _08957_ (.A(_02867_),
    .B(_02800_),
    .C(_02868_),
    .Y(_02869_));
 sky130_fd_sc_hd__nand3_1 _08958_ (.A(_02866_),
    .B(_02869_),
    .C(_00581_),
    .Y(_02870_));
 sky130_fd_sc_hd__o21ai_2 _08959_ (.A1(_00580_),
    .A2(_00671_),
    .B1(_02539_),
    .Y(_02871_));
 sky130_fd_sc_hd__inv_2 _08960_ (.A(_02871_),
    .Y(_02872_));
 sky130_fd_sc_hd__nand2_1 _08961_ (.A(_02870_),
    .B(_02872_),
    .Y(_02873_));
 sky130_fd_sc_hd__clkbuf_4 _08962_ (.A(_00006_),
    .X(_02874_));
 sky130_fd_sc_hd__nor2_1 _08963_ (.A(_02874_),
    .B(_02226_),
    .Y(_02875_));
 sky130_fd_sc_hd__nand2_1 _08964_ (.A(_02561_),
    .B(\Oset[1][3] ),
    .Y(_02876_));
 sky130_fd_sc_hd__nand2_1 _08965_ (.A(_02876_),
    .B(_02534_),
    .Y(_02877_));
 sky130_fd_sc_hd__nand2_1 _08966_ (.A(_02522_),
    .B(\Oset[2][3] ),
    .Y(_02878_));
 sky130_fd_sc_hd__nand2_1 _08967_ (.A(_02874_),
    .B(\Oset[3][3] ),
    .Y(_02879_));
 sky130_fd_sc_hd__nand3_1 _08968_ (.A(_02878_),
    .B(_02727_),
    .C(_02879_),
    .Y(_02880_));
 sky130_fd_sc_hd__o21ai_4 _08969_ (.A1(_02875_),
    .A2(_02877_),
    .B1(_02880_),
    .Y(_02881_));
 sky130_fd_sc_hd__nand2_1 _08970_ (.A(_02881_),
    .B(_02551_),
    .Y(_02882_));
 sky130_fd_sc_hd__nand3_1 _08971_ (.A(_02873_),
    .B(_01154_),
    .C(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__o21ai_1 _08972_ (.A1(_01153_),
    .A2(_00671_),
    .B1(_02555_),
    .Y(_02884_));
 sky130_fd_sc_hd__inv_2 _08973_ (.A(_02884_),
    .Y(_02885_));
 sky130_fd_sc_hd__nand2_1 _08974_ (.A(_02883_),
    .B(_02885_),
    .Y(_02886_));
 sky130_fd_sc_hd__nor2_1 _08975_ (.A(_02798_),
    .B(_02234_),
    .Y(_02887_));
 sky130_fd_sc_hd__a21o_1 _08976_ (.A1(_02528_),
    .A2(\H[1][3] ),
    .B1(_02727_),
    .X(_02888_));
 sky130_fd_sc_hd__nand2_1 _08977_ (.A(_02798_),
    .B(\H[3][3] ),
    .Y(_02889_));
 sky130_fd_sc_hd__o211ai_1 _08978_ (.A1(_02798_),
    .A2(_02231_),
    .B1(_02525_),
    .C1(_02889_),
    .Y(_02890_));
 sky130_fd_sc_hd__o21ai_2 _08979_ (.A1(_02887_),
    .A2(_02888_),
    .B1(_02890_),
    .Y(_02891_));
 sky130_fd_sc_hd__a21oi_1 _08980_ (.A1(_02891_),
    .A2(_02572_),
    .B1(_00586_),
    .Y(_02892_));
 sky130_fd_sc_hd__nand2_1 _08981_ (.A(_02886_),
    .B(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__nand2_1 _08982_ (.A(_00586_),
    .B(\R2[1] ),
    .Y(_02894_));
 sky130_fd_sc_hd__nand2_4 _08983_ (.A(_02893_),
    .B(_02894_),
    .Y(_02895_));
 sky130_fd_sc_hd__nand3_1 _08984_ (.A(_02822_),
    .B(_02620_),
    .C(_02895_),
    .Y(_02896_));
 sky130_fd_sc_hd__inv_2 _08985_ (.A(_02821_),
    .Y(_02897_));
 sky130_fd_sc_hd__a21oi_1 _08986_ (.A1(_02685_),
    .A2(_02192_),
    .B1(_02897_),
    .Y(_02898_));
 sky130_fd_sc_hd__nand2_1 _08987_ (.A(_02619_),
    .B(_02895_),
    .Y(_02899_));
 sky130_fd_sc_hd__nand2_1 _08988_ (.A(_02898_),
    .B(_02899_),
    .Y(_02900_));
 sky130_fd_sc_hd__nand2_1 _08989_ (.A(_02785_),
    .B(_02734_),
    .Y(_02901_));
 sky130_fd_sc_hd__nand3_1 _08990_ (.A(_02896_),
    .B(_02900_),
    .C(_02901_),
    .Y(_02902_));
 sky130_fd_sc_hd__a21oi_1 _08991_ (.A1(_02618_),
    .A2(_02158_),
    .B1(_02897_),
    .Y(_02903_));
 sky130_fd_sc_hd__inv_2 _08992_ (.A(_02895_),
    .Y(_02904_));
 sky130_fd_sc_hd__a21oi_1 _08993_ (.A1(_02685_),
    .A2(_02192_),
    .B1(_02904_),
    .Y(_02905_));
 sky130_fd_sc_hd__nand2_1 _08994_ (.A(_02903_),
    .B(_02905_),
    .Y(_02906_));
 sky130_fd_sc_hd__inv_2 _08995_ (.A(_02901_),
    .Y(_02907_));
 sky130_fd_sc_hd__nand2_1 _08996_ (.A(_02822_),
    .B(_02899_),
    .Y(_02908_));
 sky130_fd_sc_hd__nand3_1 _08997_ (.A(_02906_),
    .B(_02907_),
    .C(_02908_),
    .Y(_02909_));
 sky130_fd_sc_hd__nand2_1 _08998_ (.A(_02902_),
    .B(_02909_),
    .Y(_02910_));
 sky130_fd_sc_hd__nor2_1 _08999_ (.A(_02736_),
    .B(_02823_),
    .Y(_02911_));
 sky130_fd_sc_hd__a21oi_2 _09000_ (.A1(_02824_),
    .A2(_02786_),
    .B1(_02911_),
    .Y(_02912_));
 sky130_fd_sc_hd__inv_2 _09001_ (.A(_02912_),
    .Y(_02913_));
 sky130_fd_sc_hd__nand2_1 _09002_ (.A(_02910_),
    .B(_02913_),
    .Y(_02914_));
 sky130_fd_sc_hd__nand3_1 _09003_ (.A(_02912_),
    .B(_02902_),
    .C(_02909_),
    .Y(_02915_));
 sky130_fd_sc_hd__nand2_1 _09004_ (.A(_02914_),
    .B(_02915_),
    .Y(_02916_));
 sky130_fd_sc_hd__nand2_1 _09005_ (.A(_02581_),
    .B(\Oset[2][3] ),
    .Y(_02917_));
 sky130_fd_sc_hd__nand2_1 _09006_ (.A(_02592_),
    .B(\Oset[3][3] ),
    .Y(_02918_));
 sky130_fd_sc_hd__nand3_1 _09007_ (.A(_02917_),
    .B(_02584_),
    .C(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__nand2_1 _09008_ (.A(_02581_),
    .B(\Oset[0][3] ),
    .Y(_02920_));
 sky130_fd_sc_hd__nand2_1 _09009_ (.A(_02585_),
    .B(\Oset[1][3] ),
    .Y(_02921_));
 sky130_fd_sc_hd__nand3_1 _09010_ (.A(_02920_),
    .B(_02590_),
    .C(_02921_),
    .Y(_02922_));
 sky130_fd_sc_hd__nand2_1 _09011_ (.A(_02919_),
    .B(_02922_),
    .Y(_02923_));
 sky130_fd_sc_hd__o21ai_1 _09012_ (.A1(_02539_),
    .A2(_02923_),
    .B1(_01153_),
    .Y(_02924_));
 sky130_fd_sc_hd__inv_2 _09013_ (.A(_02924_),
    .Y(_02925_));
 sky130_fd_sc_hd__nand2_1 _09014_ (.A(_02222_),
    .B(_02161_),
    .Y(_02926_));
 sky130_fd_sc_hd__nand2_1 _09015_ (.A(_02582_),
    .B(\Qset[2][3] ),
    .Y(_02927_));
 sky130_fd_sc_hd__nand2_1 _09016_ (.A(_02586_),
    .B(\Qset[3][3] ),
    .Y(_02928_));
 sky130_fd_sc_hd__nand3_1 _09017_ (.A(_02927_),
    .B(_02584_),
    .C(_02928_),
    .Y(_02929_));
 sky130_fd_sc_hd__nand2_1 _09018_ (.A(_02582_),
    .B(\Qset[0][3] ),
    .Y(_02930_));
 sky130_fd_sc_hd__nand2_1 _09019_ (.A(_02586_),
    .B(\Qset[1][3] ),
    .Y(_02931_));
 sky130_fd_sc_hd__nand3_1 _09020_ (.A(_02930_),
    .B(_02591_),
    .C(_02931_),
    .Y(_02932_));
 sky130_fd_sc_hd__nand2_1 _09021_ (.A(_02929_),
    .B(_02932_),
    .Y(_02933_));
 sky130_fd_sc_hd__nand2_1 _09022_ (.A(_02933_),
    .B(_00580_),
    .Y(_02934_));
 sky130_fd_sc_hd__nand3_1 _09023_ (.A(_02926_),
    .B(_02934_),
    .C(_02540_),
    .Y(_02935_));
 sky130_fd_sc_hd__nand2_1 _09024_ (.A(_02925_),
    .B(_02935_),
    .Y(_02936_));
 sky130_fd_sc_hd__a21oi_1 _09025_ (.A1(_02229_),
    .A2(_00583_),
    .B1(_02571_),
    .Y(_02937_));
 sky130_fd_sc_hd__nand2_1 _09026_ (.A(_02936_),
    .B(_02937_),
    .Y(_02938_));
 sky130_fd_sc_hd__nor2_1 _09027_ (.A(_02592_),
    .B(_02231_),
    .Y(_02939_));
 sky130_fd_sc_hd__a211o_1 _09028_ (.A1(_02592_),
    .A2(\H[3][3] ),
    .B1(_02591_),
    .C1(_02939_),
    .X(_02940_));
 sky130_fd_sc_hd__nor2_1 _09029_ (.A(_02592_),
    .B(_02234_),
    .Y(_02941_));
 sky130_fd_sc_hd__a211o_1 _09030_ (.A1(_02592_),
    .A2(\H[1][3] ),
    .B1(_00005_),
    .C1(_02941_),
    .X(_02942_));
 sky130_fd_sc_hd__nand2_1 _09031_ (.A(_02940_),
    .B(_02942_),
    .Y(_02943_));
 sky130_fd_sc_hd__inv_2 _09032_ (.A(_02943_),
    .Y(_02944_));
 sky130_fd_sc_hd__nand2_1 _09033_ (.A(_02944_),
    .B(_02572_),
    .Y(_02945_));
 sky130_fd_sc_hd__nand2_1 _09034_ (.A(_02938_),
    .B(_02945_),
    .Y(_02946_));
 sky130_fd_sc_hd__nand2_1 _09035_ (.A(_02946_),
    .B(_01552_),
    .Y(_02947_));
 sky130_fd_sc_hd__nand2_1 _09036_ (.A(_02947_),
    .B(_02237_),
    .Y(_02948_));
 sky130_fd_sc_hd__inv_2 _09037_ (.A(_02948_),
    .Y(_02949_));
 sky130_fd_sc_hd__nor2_1 _09038_ (.A(_02578_),
    .B(_02949_),
    .Y(_02950_));
 sky130_fd_sc_hd__nand2_1 _09039_ (.A(_02916_),
    .B(_02950_),
    .Y(_02951_));
 sky130_fd_sc_hd__inv_2 _09040_ (.A(_02950_),
    .Y(_02952_));
 sky130_fd_sc_hd__nand3_1 _09041_ (.A(_02914_),
    .B(_02915_),
    .C(_02952_),
    .Y(_02953_));
 sky130_fd_sc_hd__nand3_1 _09042_ (.A(_02863_),
    .B(_02951_),
    .C(_02953_),
    .Y(_02954_));
 sky130_fd_sc_hd__nand2_1 _09043_ (.A(_02951_),
    .B(_02953_),
    .Y(_02955_));
 sky130_fd_sc_hd__nand2_1 _09044_ (.A(_02955_),
    .B(_02828_),
    .Y(_02956_));
 sky130_fd_sc_hd__nand2_1 _09045_ (.A(_02954_),
    .B(_02956_),
    .Y(_02957_));
 sky130_fd_sc_hd__nand2_1 _09046_ (.A(_02895_),
    .B(_00549_),
    .Y(_02958_));
 sky130_fd_sc_hd__o21ai_1 _09047_ (.A1(_00549_),
    .A2(_02957_),
    .B1(_02958_),
    .Y(_02959_));
 sky130_fd_sc_hd__or2_1 _09048_ (.A(\Add.sub ),
    .B(_02959_),
    .X(_02960_));
 sky130_fd_sc_hd__nand2_1 _09049_ (.A(_02959_),
    .B(\Add.sub ),
    .Y(_02961_));
 sky130_fd_sc_hd__nand2_1 _09050_ (.A(_02960_),
    .B(_02961_),
    .Y(_02962_));
 sky130_fd_sc_hd__buf_6 _09051_ (.A(_02948_),
    .X(_02963_));
 sky130_fd_sc_hd__nor2_1 _09052_ (.A(_02836_),
    .B(_02231_),
    .Y(_02964_));
 sky130_fd_sc_hd__a211o_1 _09053_ (.A1(\H[3][3] ),
    .A2(_02836_),
    .B1(_02837_),
    .C1(_02964_),
    .X(_02965_));
 sky130_fd_sc_hd__nor2_1 _09054_ (.A(_02836_),
    .B(_02234_),
    .Y(_02966_));
 sky130_fd_sc_hd__a211o_1 _09055_ (.A1(\H[1][3] ),
    .A2(_02836_),
    .B1(_02840_),
    .C1(_02966_),
    .X(_02967_));
 sky130_fd_sc_hd__a21oi_1 _09056_ (.A1(\Qset[3][3] ),
    .A2(_02836_),
    .B1(_02837_),
    .Y(_02968_));
 sky130_fd_sc_hd__nand2_1 _09057_ (.A(_02632_),
    .B(\Qset[2][3] ),
    .Y(_02969_));
 sky130_fd_sc_hd__a21oi_1 _09058_ (.A1(_02632_),
    .A2(\Qset[0][3] ),
    .B1(_02840_),
    .Y(_02970_));
 sky130_fd_sc_hd__nand2_1 _09059_ (.A(\Qset[1][3] ),
    .B(_02836_),
    .Y(_02971_));
 sky130_fd_sc_hd__a221o_1 _09060_ (.A1(_02968_),
    .A2(_02969_),
    .B1(_02970_),
    .B2(_02971_),
    .C1(Oreg3),
    .X(_02972_));
 sky130_fd_sc_hd__a21oi_1 _09061_ (.A1(\Oset[3][3] ),
    .A2(_02688_),
    .B1(_02837_),
    .Y(_02973_));
 sky130_fd_sc_hd__nand2_1 _09062_ (.A(_02632_),
    .B(\Oset[2][3] ),
    .Y(_02974_));
 sky130_fd_sc_hd__a21oi_1 _09063_ (.A1(_02632_),
    .A2(\Oset[0][3] ),
    .B1(_02840_),
    .Y(_02975_));
 sky130_fd_sc_hd__nand2_1 _09064_ (.A(\Oset[1][3] ),
    .B(_02836_),
    .Y(_02976_));
 sky130_fd_sc_hd__a221o_1 _09065_ (.A1(_02973_),
    .A2(_02974_),
    .B1(_02975_),
    .B2(_02976_),
    .C1(_00646_),
    .X(_02977_));
 sky130_fd_sc_hd__a21oi_1 _09066_ (.A1(_02972_),
    .A2(_02977_),
    .B1(_01536_),
    .Y(_02978_));
 sky130_fd_sc_hd__a311o_1 _09067_ (.A1(_01536_),
    .A2(_02965_),
    .A3(_02967_),
    .B1(_00549_),
    .C1(_02978_),
    .X(_02979_));
 sky130_fd_sc_hd__o21ai_1 _09068_ (.A1(_00622_),
    .A2(_02963_),
    .B1(_02979_),
    .Y(_02980_));
 sky130_fd_sc_hd__nand2_1 _09069_ (.A(_02962_),
    .B(_02980_),
    .Y(_02981_));
 sky130_fd_sc_hd__nand3b_1 _09070_ (.A_N(_02980_),
    .B(_02960_),
    .C(_02961_),
    .Y(_02982_));
 sky130_fd_sc_hd__nand2_1 _09071_ (.A(_02859_),
    .B(_02856_),
    .Y(_02983_));
 sky130_fd_sc_hd__a21o_1 _09072_ (.A1(_02981_),
    .A2(_02982_),
    .B1(_02983_),
    .X(_02984_));
 sky130_fd_sc_hd__nand3_1 _09073_ (.A(_02983_),
    .B(_02981_),
    .C(_02982_),
    .Y(_02985_));
 sky130_fd_sc_hd__and2_2 _09074_ (.A(_02984_),
    .B(_02985_),
    .X(_02986_));
 sky130_fd_sc_hd__nor2_1 _09075_ (.A(_02653_),
    .B(_02986_),
    .Y(_02987_));
 sky130_fd_sc_hd__a211o_1 _09076_ (.A1(_00762_),
    .A2(_02654_),
    .B1(_02753_),
    .C1(_02987_),
    .X(_02988_));
 sky130_fd_sc_hd__inv_2 _09077_ (.A(_02988_),
    .Y(_00247_));
 sky130_fd_sc_hd__nand2_1 _09078_ (.A(_02247_),
    .B(_02161_),
    .Y(_02989_));
 sky130_fd_sc_hd__nand2_1 _09079_ (.A(_02582_),
    .B(\Qset[2][4] ),
    .Y(_02990_));
 sky130_fd_sc_hd__buf_4 _09080_ (.A(_02584_),
    .X(_02991_));
 sky130_fd_sc_hd__buf_6 _09081_ (.A(_02586_),
    .X(_02992_));
 sky130_fd_sc_hd__nand2_1 _09082_ (.A(_02992_),
    .B(\Qset[3][4] ),
    .Y(_02993_));
 sky130_fd_sc_hd__nand3_1 _09083_ (.A(_02990_),
    .B(_02991_),
    .C(_02993_),
    .Y(_02994_));
 sky130_fd_sc_hd__nand2_1 _09084_ (.A(_02582_),
    .B(\Qset[0][4] ),
    .Y(_02995_));
 sky130_fd_sc_hd__nand2_1 _09085_ (.A(_02992_),
    .B(\Qset[1][4] ),
    .Y(_02996_));
 sky130_fd_sc_hd__nand3_1 _09086_ (.A(_02995_),
    .B(_02591_),
    .C(_02996_),
    .Y(_02997_));
 sky130_fd_sc_hd__nand2_1 _09087_ (.A(_02994_),
    .B(_02997_),
    .Y(_02998_));
 sky130_fd_sc_hd__nand2_1 _09088_ (.A(_02998_),
    .B(_00581_),
    .Y(_02999_));
 sky130_fd_sc_hd__nand3_1 _09089_ (.A(_02989_),
    .B(_02999_),
    .C(_02540_),
    .Y(_03000_));
 sky130_fd_sc_hd__buf_6 _09090_ (.A(_02611_),
    .X(_03001_));
 sky130_fd_sc_hd__nand2_1 _09091_ (.A(_03001_),
    .B(\Oset[3][4] ),
    .Y(_03002_));
 sky130_fd_sc_hd__o211ai_1 _09092_ (.A1(_03001_),
    .A2(_02249_),
    .B1(_02991_),
    .C1(_03002_),
    .Y(_03003_));
 sky130_fd_sc_hd__buf_6 _09093_ (.A(_02591_),
    .X(_03004_));
 sky130_fd_sc_hd__nand2_1 _09094_ (.A(_03001_),
    .B(\Oset[1][4] ),
    .Y(_03005_));
 sky130_fd_sc_hd__o211ai_1 _09095_ (.A1(_02992_),
    .A2(_02253_),
    .B1(_03004_),
    .C1(_03005_),
    .Y(_03006_));
 sky130_fd_sc_hd__nand3_1 _09096_ (.A(_03003_),
    .B(_03006_),
    .C(_02551_),
    .Y(_03007_));
 sky130_fd_sc_hd__nand3_1 _09097_ (.A(_03000_),
    .B(_01154_),
    .C(_03007_),
    .Y(_03008_));
 sky130_fd_sc_hd__a21oi_1 _09098_ (.A1(_02257_),
    .A2(_00583_),
    .B1(_02572_),
    .Y(_03009_));
 sky130_fd_sc_hd__nand2_1 _09099_ (.A(_03008_),
    .B(_03009_),
    .Y(_03010_));
 sky130_fd_sc_hd__nor2_1 _09100_ (.A(\H[3][4] ),
    .B(_02582_),
    .Y(_03011_));
 sky130_fd_sc_hd__o21ai_1 _09101_ (.A1(_02611_),
    .A2(\H[2][4] ),
    .B1(_02584_),
    .Y(_03012_));
 sky130_fd_sc_hd__nor2_1 _09102_ (.A(_02611_),
    .B(\H[0][4] ),
    .Y(_03013_));
 sky130_fd_sc_hd__o21ai_1 _09103_ (.A1(\H[1][4] ),
    .A2(_02582_),
    .B1(_02591_),
    .Y(_03014_));
 sky130_fd_sc_hd__o22a_1 _09104_ (.A1(_03011_),
    .A2(_03012_),
    .B1(_03013_),
    .B2(_03014_),
    .X(_03015_));
 sky130_fd_sc_hd__or2_1 _09105_ (.A(_02556_),
    .B(_03015_),
    .X(_03016_));
 sky130_fd_sc_hd__nand2_1 _09106_ (.A(_03010_),
    .B(_03016_),
    .Y(_03017_));
 sky130_fd_sc_hd__nand2_2 _09107_ (.A(_03017_),
    .B(_01552_),
    .Y(_03018_));
 sky130_fd_sc_hd__nand2_2 _09108_ (.A(_03018_),
    .B(_02264_),
    .Y(_03019_));
 sky130_fd_sc_hd__buf_6 _09109_ (.A(_03019_),
    .X(_03020_));
 sky130_fd_sc_hd__buf_2 _09110_ (.A(_02632_),
    .X(_03021_));
 sky130_fd_sc_hd__clkbuf_4 _09111_ (.A(_03021_),
    .X(_03022_));
 sky130_fd_sc_hd__clkbuf_4 _09112_ (.A(_03022_),
    .X(_03023_));
 sky130_fd_sc_hd__buf_2 _09113_ (.A(_02836_),
    .X(_03024_));
 sky130_fd_sc_hd__clkbuf_4 _09114_ (.A(_03024_),
    .X(_03025_));
 sky130_fd_sc_hd__buf_2 _09115_ (.A(_02837_),
    .X(_03026_));
 sky130_fd_sc_hd__clkbuf_4 _09116_ (.A(_03026_),
    .X(_03027_));
 sky130_fd_sc_hd__a21o_1 _09117_ (.A1(\H[3][4] ),
    .A2(_03025_),
    .B1(_03027_),
    .X(_03028_));
 sky130_fd_sc_hd__a21o_1 _09118_ (.A1(\H[2][4] ),
    .A2(_03023_),
    .B1(_03028_),
    .X(_03029_));
 sky130_fd_sc_hd__a21o_1 _09119_ (.A1(\H[1][4] ),
    .A2(_03025_),
    .B1(_02840_),
    .X(_03030_));
 sky130_fd_sc_hd__a21o_1 _09120_ (.A1(\H[0][4] ),
    .A2(_03023_),
    .B1(_03030_),
    .X(_03031_));
 sky130_fd_sc_hd__nand2_1 _09121_ (.A(_03022_),
    .B(\Qset[0][4] ),
    .Y(_03032_));
 sky130_fd_sc_hd__buf_2 _09122_ (.A(_03024_),
    .X(_03033_));
 sky130_fd_sc_hd__nand2_1 _09123_ (.A(\Qset[1][4] ),
    .B(_03033_),
    .Y(_03034_));
 sky130_fd_sc_hd__a21oi_1 _09124_ (.A1(\Qset[3][4] ),
    .A2(_03025_),
    .B1(_03027_),
    .Y(_03035_));
 sky130_fd_sc_hd__nand2_1 _09125_ (.A(_03022_),
    .B(\Qset[2][4] ),
    .Y(_03036_));
 sky130_fd_sc_hd__a32o_1 _09126_ (.A1(_03032_),
    .A2(_03034_),
    .A3(_03027_),
    .B1(_03035_),
    .B2(_03036_),
    .X(_03037_));
 sky130_fd_sc_hd__nand2_1 _09127_ (.A(_03022_),
    .B(\Oset[0][4] ),
    .Y(_03038_));
 sky130_fd_sc_hd__nand2_1 _09128_ (.A(\Oset[1][4] ),
    .B(_03033_),
    .Y(_03039_));
 sky130_fd_sc_hd__a21oi_1 _09129_ (.A1(\Oset[3][4] ),
    .A2(_03025_),
    .B1(_03027_),
    .Y(_03040_));
 sky130_fd_sc_hd__nand2_1 _09130_ (.A(_03022_),
    .B(\Oset[2][4] ),
    .Y(_03041_));
 sky130_fd_sc_hd__a32o_1 _09131_ (.A1(_03038_),
    .A2(_03039_),
    .A3(_03027_),
    .B1(_03040_),
    .B2(_03041_),
    .X(_03042_));
 sky130_fd_sc_hd__mux2_1 _09132_ (.A0(_03037_),
    .A1(_03042_),
    .S(_00621_),
    .X(_03043_));
 sky130_fd_sc_hd__nor2_1 _09133_ (.A(_01537_),
    .B(_03043_),
    .Y(_03044_));
 sky130_fd_sc_hd__a311o_2 _09134_ (.A1(_01537_),
    .A2(_03029_),
    .A3(_03031_),
    .B1(_00556_),
    .C1(_03044_),
    .X(_03045_));
 sky130_fd_sc_hd__o21ai_2 _09135_ (.A1(_00624_),
    .A2(_03020_),
    .B1(_03045_),
    .Y(_03046_));
 sky130_fd_sc_hd__nor2_1 _09136_ (.A(_00583_),
    .B(_02551_),
    .Y(_03047_));
 sky130_fd_sc_hd__inv_2 _09137_ (.A(_03047_),
    .Y(_03048_));
 sky130_fd_sc_hd__nor2_4 _09138_ (.A(\shift.H ),
    .B(_02571_),
    .Y(_03049_));
 sky130_fd_sc_hd__inv_6 _09139_ (.A(_03049_),
    .Y(_03050_));
 sky130_fd_sc_hd__nor2_2 _09140_ (.A(_03048_),
    .B(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hd__nor2_1 _09141_ (.A(_03051_),
    .B(_02738_),
    .Y(_03052_));
 sky130_fd_sc_hd__nor2_1 _09142_ (.A(_02874_),
    .B(_02312_),
    .Y(_03053_));
 sky130_fd_sc_hd__a211o_1 _09143_ (.A1(_02528_),
    .A2(\Qset[3][7] ),
    .B1(_02534_),
    .C1(_03053_),
    .X(_03054_));
 sky130_fd_sc_hd__nor2_1 _09144_ (.A(_02561_),
    .B(_02315_),
    .Y(_03055_));
 sky130_fd_sc_hd__a211o_1 _09145_ (.A1(_02528_),
    .A2(\Qset[1][7] ),
    .B1(_02727_),
    .C1(_03055_),
    .X(_03056_));
 sky130_fd_sc_hd__nand3_1 _09146_ (.A(_03054_),
    .B(_03056_),
    .C(_00581_),
    .Y(_03057_));
 sky130_fd_sc_hd__nand2_1 _09147_ (.A(_03057_),
    .B(_02872_),
    .Y(_03058_));
 sky130_fd_sc_hd__nor2_1 _09148_ (.A(_02561_),
    .B(_02320_),
    .Y(_03059_));
 sky130_fd_sc_hd__a211o_1 _09149_ (.A1(_02874_),
    .A2(\Oset[3][7] ),
    .B1(_02534_),
    .C1(_03059_),
    .X(_03060_));
 sky130_fd_sc_hd__nor2_1 _09150_ (.A(_02561_),
    .B(_02323_),
    .Y(_03061_));
 sky130_fd_sc_hd__a211o_1 _09151_ (.A1(_02874_),
    .A2(\Oset[1][7] ),
    .B1(_02727_),
    .C1(_03061_),
    .X(_03062_));
 sky130_fd_sc_hd__nand2_2 _09152_ (.A(_03060_),
    .B(_03062_),
    .Y(_03063_));
 sky130_fd_sc_hd__nand2_1 _09153_ (.A(_03063_),
    .B(_02552_),
    .Y(_03064_));
 sky130_fd_sc_hd__nand3_1 _09154_ (.A(_03058_),
    .B(_01154_),
    .C(_03064_),
    .Y(_03065_));
 sky130_fd_sc_hd__o21ai_2 _09155_ (.A1(_01154_),
    .A2(_01990_),
    .B1(_02555_),
    .Y(_03066_));
 sky130_fd_sc_hd__inv_2 _09156_ (.A(_03066_),
    .Y(_03067_));
 sky130_fd_sc_hd__nand2_1 _09157_ (.A(_03065_),
    .B(_03067_),
    .Y(_03068_));
 sky130_fd_sc_hd__or2_1 _09158_ (.A(_02874_),
    .B(\H[0][7] ),
    .X(_03069_));
 sky130_fd_sc_hd__o21a_1 _09159_ (.A1(\H[1][7] ),
    .A2(_02522_),
    .B1(_02800_),
    .X(_03070_));
 sky130_fd_sc_hd__mux2_1 _09160_ (.A0(\H[2][7] ),
    .A1(\H[3][7] ),
    .S(_02561_),
    .X(_03071_));
 sky130_fd_sc_hd__a22oi_4 _09161_ (.A1(_03069_),
    .A2(_03070_),
    .B1(_03071_),
    .B2(_02526_),
    .Y(_03072_));
 sky130_fd_sc_hd__a21oi_1 _09162_ (.A1(_03072_),
    .A2(_02572_),
    .B1(_00586_),
    .Y(_03073_));
 sky130_fd_sc_hd__nand2_1 _09163_ (.A(_03068_),
    .B(_03073_),
    .Y(_03074_));
 sky130_fd_sc_hd__nand2_1 _09164_ (.A(_00587_),
    .B(\im_reg[7] ),
    .Y(_03075_));
 sky130_fd_sc_hd__nand2_4 _09165_ (.A(_03074_),
    .B(_03075_),
    .Y(_03076_));
 sky130_fd_sc_hd__nand2_1 _09166_ (.A(_03052_),
    .B(_03076_),
    .Y(_03077_));
 sky130_fd_sc_hd__inv_2 _09167_ (.A(_03077_),
    .Y(_03078_));
 sky130_fd_sc_hd__inv_2 _09168_ (.A(_03051_),
    .Y(_03079_));
 sky130_fd_sc_hd__and2_1 _09169_ (.A(_02619_),
    .B(_03079_),
    .X(_03080_));
 sky130_fd_sc_hd__nor2_1 _09170_ (.A(_02528_),
    .B(_02292_),
    .Y(_03081_));
 sky130_fd_sc_hd__a211o_1 _09171_ (.A1(_02544_),
    .A2(\Qset[1][6] ),
    .B1(_02727_),
    .C1(_03081_),
    .X(_03082_));
 sky130_fd_sc_hd__nor2_1 _09172_ (.A(_02528_),
    .B(_02289_),
    .Y(_03083_));
 sky130_fd_sc_hd__a211o_1 _09173_ (.A1(_02544_),
    .A2(\Qset[3][6] ),
    .B1(_02800_),
    .C1(_03083_),
    .X(_03084_));
 sky130_fd_sc_hd__nand3_1 _09174_ (.A(_03082_),
    .B(_03084_),
    .C(_00581_),
    .Y(_03085_));
 sky130_fd_sc_hd__nand2_1 _09175_ (.A(_03085_),
    .B(_02796_),
    .Y(_03086_));
 sky130_fd_sc_hd__nor2_1 _09176_ (.A(_02874_),
    .B(_02296_),
    .Y(_03087_));
 sky130_fd_sc_hd__a211o_1 _09177_ (.A1(_02544_),
    .A2(\Oset[3][6] ),
    .B1(_02534_),
    .C1(_03087_),
    .X(_03088_));
 sky130_fd_sc_hd__nor2_1 _09178_ (.A(_02874_),
    .B(_02299_),
    .Y(_03089_));
 sky130_fd_sc_hd__a211o_1 _09179_ (.A1(_02544_),
    .A2(\Oset[1][6] ),
    .B1(_02727_),
    .C1(_03089_),
    .X(_03090_));
 sky130_fd_sc_hd__nand2_2 _09180_ (.A(_03088_),
    .B(_03090_),
    .Y(_03091_));
 sky130_fd_sc_hd__nand2_1 _09181_ (.A(_03091_),
    .B(_02552_),
    .Y(_03092_));
 sky130_fd_sc_hd__nand3_1 _09182_ (.A(_03086_),
    .B(_01155_),
    .C(_03092_),
    .Y(_03093_));
 sky130_fd_sc_hd__inv_2 _09183_ (.A(\im_reg[6] ),
    .Y(_03094_));
 sky130_fd_sc_hd__o21ai_2 _09184_ (.A1(_01154_),
    .A2(_03094_),
    .B1(_02555_),
    .Y(_03095_));
 sky130_fd_sc_hd__inv_2 _09185_ (.A(_03095_),
    .Y(_03096_));
 sky130_fd_sc_hd__nand2_1 _09186_ (.A(_03093_),
    .B(_03096_),
    .Y(_03097_));
 sky130_fd_sc_hd__nand2_1 _09187_ (.A(_02787_),
    .B(\H[0][6] ),
    .Y(_03098_));
 sky130_fd_sc_hd__nand2_1 _09188_ (.A(_02562_),
    .B(\H[1][6] ),
    .Y(_03099_));
 sky130_fd_sc_hd__a21o_1 _09189_ (.A1(_02874_),
    .A2(\H[3][6] ),
    .B1(_02534_),
    .X(_03100_));
 sky130_fd_sc_hd__a21oi_1 _09190_ (.A1(_02787_),
    .A2(\H[2][6] ),
    .B1(_03100_),
    .Y(_03101_));
 sky130_fd_sc_hd__a31o_2 _09191_ (.A1(_02535_),
    .A2(_03098_),
    .A3(_03099_),
    .B1(_03101_),
    .X(_03102_));
 sky130_fd_sc_hd__a21oi_1 _09192_ (.A1(_03102_),
    .A2(_02572_),
    .B1(_00586_),
    .Y(_03103_));
 sky130_fd_sc_hd__nand2_1 _09193_ (.A(_03097_),
    .B(_03103_),
    .Y(_03104_));
 sky130_fd_sc_hd__nand2_1 _09194_ (.A(_00587_),
    .B(\im_reg[6] ),
    .Y(_03105_));
 sky130_fd_sc_hd__nand2_2 _09195_ (.A(_03104_),
    .B(_03105_),
    .Y(_03106_));
 sky130_fd_sc_hd__nand2_1 _09196_ (.A(_03080_),
    .B(_03106_),
    .Y(_03107_));
 sky130_fd_sc_hd__inv_2 _09197_ (.A(_03107_),
    .Y(_03108_));
 sky130_fd_sc_hd__nand2_1 _09198_ (.A(_03078_),
    .B(_03108_),
    .Y(_03109_));
 sky130_fd_sc_hd__clkbuf_4 _09199_ (.A(_03106_),
    .X(_03110_));
 sky130_fd_sc_hd__nand2_1 _09200_ (.A(_03052_),
    .B(_03110_),
    .Y(_03111_));
 sky130_fd_sc_hd__nand2_1 _09201_ (.A(_03080_),
    .B(_03076_),
    .Y(_03112_));
 sky130_fd_sc_hd__nand2_1 _09202_ (.A(_03111_),
    .B(_03112_),
    .Y(_03113_));
 sky130_fd_sc_hd__nand2_1 _09203_ (.A(_03109_),
    .B(_03113_),
    .Y(_03114_));
 sky130_fd_sc_hd__inv_2 _09204_ (.A(_02784_),
    .Y(_03115_));
 sky130_fd_sc_hd__nor2_1 _09205_ (.A(_03051_),
    .B(_03115_),
    .Y(_03116_));
 sky130_fd_sc_hd__nor2_1 _09206_ (.A(_02529_),
    .B(_02277_),
    .Y(_03117_));
 sky130_fd_sc_hd__nand2_1 _09207_ (.A(_02544_),
    .B(\Oset[1][5] ),
    .Y(_03118_));
 sky130_fd_sc_hd__inv_2 _09208_ (.A(_03118_),
    .Y(_03119_));
 sky130_fd_sc_hd__nor2_1 _09209_ (.A(_02798_),
    .B(_02274_),
    .Y(_03120_));
 sky130_fd_sc_hd__a211o_1 _09210_ (.A1(_02562_),
    .A2(\Oset[3][5] ),
    .B1(_02800_),
    .C1(_03120_),
    .X(_03121_));
 sky130_fd_sc_hd__o31ai_4 _09211_ (.A1(_02525_),
    .A2(_03117_),
    .A3(_03119_),
    .B1(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__nand2_1 _09212_ (.A(_03122_),
    .B(_02552_),
    .Y(_03123_));
 sky130_fd_sc_hd__a21o_1 _09213_ (.A1(_02528_),
    .A2(\Qset[3][5] ),
    .B1(_02534_),
    .X(_03124_));
 sky130_fd_sc_hd__a21o_1 _09214_ (.A1(_02523_),
    .A2(\Qset[2][5] ),
    .B1(_03124_),
    .X(_03125_));
 sky130_fd_sc_hd__a21o_1 _09215_ (.A1(_02528_),
    .A2(\Qset[1][5] ),
    .B1(_02727_),
    .X(_03126_));
 sky130_fd_sc_hd__a21o_1 _09216_ (.A1(_02787_),
    .A2(\Qset[0][5] ),
    .B1(_03126_),
    .X(_03127_));
 sky130_fd_sc_hd__nand2_2 _09217_ (.A(_03125_),
    .B(_03127_),
    .Y(_03128_));
 sky130_fd_sc_hd__o21ai_1 _09218_ (.A1(_02161_),
    .A2(_03128_),
    .B1(_02713_),
    .Y(_03129_));
 sky130_fd_sc_hd__nand3_1 _09219_ (.A(_03123_),
    .B(_03129_),
    .C(_01155_),
    .Y(_03130_));
 sky130_fd_sc_hd__nand2_1 _09220_ (.A(_00583_),
    .B(\R1[1] ),
    .Y(_03131_));
 sky130_fd_sc_hd__nand2_1 _09221_ (.A(_02556_),
    .B(_03131_),
    .Y(_03132_));
 sky130_fd_sc_hd__inv_2 _09222_ (.A(_03132_),
    .Y(_03133_));
 sky130_fd_sc_hd__nand2_1 _09223_ (.A(_03130_),
    .B(_03133_),
    .Y(_03134_));
 sky130_fd_sc_hd__buf_4 _09224_ (.A(_02800_),
    .X(_03135_));
 sky130_fd_sc_hd__buf_4 _09225_ (.A(_02787_),
    .X(_03136_));
 sky130_fd_sc_hd__nand2_1 _09226_ (.A(_03136_),
    .B(\H[0][5] ),
    .Y(_03137_));
 sky130_fd_sc_hd__nand2_1 _09227_ (.A(_02545_),
    .B(\H[1][5] ),
    .Y(_03138_));
 sky130_fd_sc_hd__a21o_1 _09228_ (.A1(_02798_),
    .A2(\H[3][5] ),
    .B1(_02800_),
    .X(_03139_));
 sky130_fd_sc_hd__a21oi_1 _09229_ (.A1(_03136_),
    .A2(\H[2][5] ),
    .B1(_03139_),
    .Y(_03140_));
 sky130_fd_sc_hd__a31o_2 _09230_ (.A1(_03135_),
    .A2(_03137_),
    .A3(_03138_),
    .B1(_03140_),
    .X(_03141_));
 sky130_fd_sc_hd__a21oi_1 _09231_ (.A1(_03141_),
    .A2(_02573_),
    .B1(_00587_),
    .Y(_03142_));
 sky130_fd_sc_hd__nand2_1 _09232_ (.A(_03134_),
    .B(_03142_),
    .Y(_03143_));
 sky130_fd_sc_hd__nand2_1 _09233_ (.A(_00587_),
    .B(\R1[1] ),
    .Y(_03144_));
 sky130_fd_sc_hd__nand2_4 _09234_ (.A(_03143_),
    .B(_03144_),
    .Y(_03145_));
 sky130_fd_sc_hd__nand2_1 _09235_ (.A(_03116_),
    .B(_03145_),
    .Y(_03146_));
 sky130_fd_sc_hd__inv_2 _09236_ (.A(_03146_),
    .Y(_03147_));
 sky130_fd_sc_hd__nand2b_1 _09237_ (.A_N(_03114_),
    .B(_03147_),
    .Y(_03148_));
 sky130_fd_sc_hd__nand2_1 _09238_ (.A(_03114_),
    .B(_03146_),
    .Y(_03149_));
 sky130_fd_sc_hd__nand2_1 _09239_ (.A(_03148_),
    .B(_03149_),
    .Y(_03150_));
 sky130_fd_sc_hd__mux2_1 _09240_ (.A0(\H[0][4] ),
    .A1(\H[1][4] ),
    .S(_02562_),
    .X(_03151_));
 sky130_fd_sc_hd__buf_4 _09241_ (.A(_02523_),
    .X(_03152_));
 sky130_fd_sc_hd__nand2_1 _09242_ (.A(_03152_),
    .B(\H[2][4] ),
    .Y(_03153_));
 sky130_fd_sc_hd__a21oi_1 _09243_ (.A1(_02567_),
    .A2(\H[3][4] ),
    .B1(_03135_),
    .Y(_03154_));
 sky130_fd_sc_hd__a2bb2o_2 _09244_ (.A1_N(_02560_),
    .A2_N(_03151_),
    .B1(_03153_),
    .B2(_03154_),
    .X(_03155_));
 sky130_fd_sc_hd__a21oi_1 _09245_ (.A1(_03155_),
    .A2(_02573_),
    .B1(_00588_),
    .Y(_03156_));
 sky130_fd_sc_hd__buf_4 _09246_ (.A(_02798_),
    .X(_03157_));
 sky130_fd_sc_hd__and2b_1 _09247_ (.A_N(_02544_),
    .B(\Qset[0][4] ),
    .X(_03158_));
 sky130_fd_sc_hd__a211o_1 _09248_ (.A1(_03157_),
    .A2(\Qset[1][4] ),
    .B1(_02526_),
    .C1(_03158_),
    .X(_03159_));
 sky130_fd_sc_hd__a21o_1 _09249_ (.A1(_02562_),
    .A2(\Qset[3][4] ),
    .B1(_02800_),
    .X(_03160_));
 sky130_fd_sc_hd__a21o_1 _09250_ (.A1(_03136_),
    .A2(\Qset[2][4] ),
    .B1(_03160_),
    .X(_03161_));
 sky130_fd_sc_hd__nand2_1 _09251_ (.A(_03159_),
    .B(_03161_),
    .Y(_03162_));
 sky130_fd_sc_hd__o21ai_1 _09252_ (.A1(_02162_),
    .A2(_03162_),
    .B1(_02542_),
    .Y(_03163_));
 sky130_fd_sc_hd__nor2_1 _09253_ (.A(_02565_),
    .B(_02253_),
    .Y(_03164_));
 sky130_fd_sc_hd__nand2_1 _09254_ (.A(_02562_),
    .B(\Oset[1][4] ),
    .Y(_03165_));
 sky130_fd_sc_hd__inv_2 _09255_ (.A(_03165_),
    .Y(_03166_));
 sky130_fd_sc_hd__nor2_1 _09256_ (.A(_02545_),
    .B(_02249_),
    .Y(_03167_));
 sky130_fd_sc_hd__a211o_1 _09257_ (.A1(_03157_),
    .A2(\Oset[3][4] ),
    .B1(_02535_),
    .C1(_03167_),
    .X(_03168_));
 sky130_fd_sc_hd__o31ai_4 _09258_ (.A1(_02560_),
    .A2(_03164_),
    .A3(_03166_),
    .B1(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hd__nand2_1 _09259_ (.A(_03169_),
    .B(_02552_),
    .Y(_03170_));
 sky130_fd_sc_hd__nand3_1 _09260_ (.A(_03163_),
    .B(_01155_),
    .C(_03170_),
    .Y(_03171_));
 sky130_fd_sc_hd__nand2_1 _09261_ (.A(\R1[0] ),
    .B(_00584_),
    .Y(_03172_));
 sky130_fd_sc_hd__nand3_1 _09262_ (.A(_03171_),
    .B(_02556_),
    .C(_03172_),
    .Y(_03173_));
 sky130_fd_sc_hd__nand2_1 _09263_ (.A(_03156_),
    .B(_03173_),
    .Y(_03174_));
 sky130_fd_sc_hd__nand2_1 _09264_ (.A(_00498_),
    .B(_00588_),
    .Y(_03175_));
 sky130_fd_sc_hd__nand2_2 _09265_ (.A(_03174_),
    .B(_03175_),
    .Y(_03176_));
 sky130_fd_sc_hd__nand2_1 _09266_ (.A(_03176_),
    .B(_03116_),
    .Y(_03177_));
 sky130_fd_sc_hd__inv_2 _09267_ (.A(_03177_),
    .Y(_03178_));
 sky130_fd_sc_hd__nand2_1 _09268_ (.A(_03052_),
    .B(_03145_),
    .Y(_03179_));
 sky130_fd_sc_hd__nand2_1 _09269_ (.A(_03179_),
    .B(_03107_),
    .Y(_03180_));
 sky130_fd_sc_hd__nor2_1 _09270_ (.A(_03107_),
    .B(_03179_),
    .Y(_03181_));
 sky130_fd_sc_hd__a21oi_1 _09271_ (.A1(_03178_),
    .A2(_03180_),
    .B1(_03181_),
    .Y(_03182_));
 sky130_fd_sc_hd__nand2_1 _09272_ (.A(_03150_),
    .B(_03182_),
    .Y(_03183_));
 sky130_fd_sc_hd__nor2_1 _09273_ (.A(_03051_),
    .B(_02949_),
    .Y(_03184_));
 sky130_fd_sc_hd__nand2_1 _09274_ (.A(_03176_),
    .B(_03184_),
    .Y(_03185_));
 sky130_fd_sc_hd__inv_2 _09275_ (.A(_03185_),
    .Y(_03186_));
 sky130_fd_sc_hd__nand3b_2 _09276_ (.A_N(_03182_),
    .B(_03148_),
    .C(_03149_),
    .Y(_03187_));
 sky130_fd_sc_hd__inv_2 _09277_ (.A(_03187_),
    .Y(_03188_));
 sky130_fd_sc_hd__a21oi_1 _09278_ (.A1(_03183_),
    .A2(_03186_),
    .B1(_03188_),
    .Y(_03189_));
 sky130_fd_sc_hd__nand2_1 _09279_ (.A(_03116_),
    .B(_03106_),
    .Y(_03190_));
 sky130_fd_sc_hd__nor2_1 _09280_ (.A(_03077_),
    .B(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hd__nand2_1 _09281_ (.A(_03077_),
    .B(_03190_),
    .Y(_03192_));
 sky130_fd_sc_hd__inv_2 _09282_ (.A(_03192_),
    .Y(_03193_));
 sky130_fd_sc_hd__nand2_1 _09283_ (.A(_03184_),
    .B(_03145_),
    .Y(_03194_));
 sky130_fd_sc_hd__o21ai_1 _09284_ (.A1(_03191_),
    .A2(_03193_),
    .B1(_03194_),
    .Y(_03195_));
 sky130_fd_sc_hd__nor2_1 _09285_ (.A(_03191_),
    .B(_03193_),
    .Y(_03196_));
 sky130_fd_sc_hd__inv_2 _09286_ (.A(_03194_),
    .Y(_03197_));
 sky130_fd_sc_hd__nand2_1 _09287_ (.A(_03196_),
    .B(_03197_),
    .Y(_03198_));
 sky130_fd_sc_hd__nand2_1 _09288_ (.A(_03195_),
    .B(_03198_),
    .Y(_03199_));
 sky130_fd_sc_hd__inv_2 _09289_ (.A(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__o21a_1 _09290_ (.A1(_03146_),
    .A2(_03114_),
    .B1(_03109_),
    .X(_03201_));
 sky130_fd_sc_hd__nand2_1 _09291_ (.A(_03200_),
    .B(_03201_),
    .Y(_03202_));
 sky130_fd_sc_hd__nand2_1 _09292_ (.A(_03148_),
    .B(_03109_),
    .Y(_03203_));
 sky130_fd_sc_hd__nand2_1 _09293_ (.A(_03203_),
    .B(_03199_),
    .Y(_03204_));
 sky130_fd_sc_hd__inv_2 _09294_ (.A(_03020_),
    .Y(_03205_));
 sky130_fd_sc_hd__inv_2 _09295_ (.A(_03176_),
    .Y(_03206_));
 sky130_fd_sc_hd__nor2_1 _09296_ (.A(_03205_),
    .B(_03206_),
    .Y(_03207_));
 sky130_fd_sc_hd__inv_2 _09297_ (.A(_03207_),
    .Y(_03208_));
 sky130_fd_sc_hd__nand3_1 _09298_ (.A(_03202_),
    .B(_03204_),
    .C(_03208_),
    .Y(_03209_));
 sky130_fd_sc_hd__nand2_1 _09299_ (.A(_03200_),
    .B(_03203_),
    .Y(_03210_));
 sky130_fd_sc_hd__nand2_1 _09300_ (.A(_03201_),
    .B(_03199_),
    .Y(_03211_));
 sky130_fd_sc_hd__nand3_1 _09301_ (.A(_03210_),
    .B(_03211_),
    .C(_03207_),
    .Y(_03212_));
 sky130_fd_sc_hd__nand2_1 _09302_ (.A(_03209_),
    .B(_03212_),
    .Y(_03213_));
 sky130_fd_sc_hd__nor2_1 _09303_ (.A(_03189_),
    .B(_03213_),
    .Y(_03214_));
 sky130_fd_sc_hd__nand2_1 _09304_ (.A(_03213_),
    .B(_03189_),
    .Y(_03215_));
 sky130_fd_sc_hd__inv_2 _09305_ (.A(_03215_),
    .Y(_03216_));
 sky130_fd_sc_hd__nand2_1 _09306_ (.A(_03187_),
    .B(_03183_),
    .Y(_03217_));
 sky130_fd_sc_hd__nand2_1 _09307_ (.A(_03217_),
    .B(_03185_),
    .Y(_03218_));
 sky130_fd_sc_hd__nand3_1 _09308_ (.A(_03187_),
    .B(_03183_),
    .C(_03186_),
    .Y(_03219_));
 sky130_fd_sc_hd__nand2_1 _09309_ (.A(_03145_),
    .B(_03080_),
    .Y(_03220_));
 sky130_fd_sc_hd__o21ai_1 _09310_ (.A1(_03220_),
    .A2(_03111_),
    .B1(_03180_),
    .Y(_03221_));
 sky130_fd_sc_hd__xor2_1 _09311_ (.A(_03178_),
    .B(_03221_),
    .X(_03222_));
 sky130_fd_sc_hd__inv_2 _09312_ (.A(_03222_),
    .Y(_03223_));
 sky130_fd_sc_hd__nand2_1 _09313_ (.A(_03176_),
    .B(_03080_),
    .Y(_03224_));
 sky130_fd_sc_hd__nor2_1 _09314_ (.A(_03179_),
    .B(_03224_),
    .Y(_03225_));
 sky130_fd_sc_hd__nand2_1 _09315_ (.A(_03223_),
    .B(_03225_),
    .Y(_03226_));
 sky130_fd_sc_hd__inv_2 _09316_ (.A(_03226_),
    .Y(_03227_));
 sky130_fd_sc_hd__nand3_2 _09317_ (.A(_03218_),
    .B(_03219_),
    .C(_03227_),
    .Y(_03228_));
 sky130_fd_sc_hd__o21ai_1 _09318_ (.A1(_03214_),
    .A2(_03216_),
    .B1(_03228_),
    .Y(_03229_));
 sky130_fd_sc_hd__nor2_1 _09319_ (.A(_03214_),
    .B(_03216_),
    .Y(_03230_));
 sky130_fd_sc_hd__inv_2 _09320_ (.A(_03228_),
    .Y(_03231_));
 sky130_fd_sc_hd__nand2_1 _09321_ (.A(_03230_),
    .B(_03231_),
    .Y(_03232_));
 sky130_fd_sc_hd__clkbuf_4 _09322_ (.A(_03051_),
    .X(_03233_));
 sky130_fd_sc_hd__nand3_1 _09323_ (.A(_03229_),
    .B(_03232_),
    .C(_03233_),
    .Y(_03234_));
 sky130_fd_sc_hd__nand2_1 _09324_ (.A(_02910_),
    .B(_02912_),
    .Y(_03235_));
 sky130_fd_sc_hd__nor2_1 _09325_ (.A(_02912_),
    .B(_02910_),
    .Y(_03236_));
 sky130_fd_sc_hd__a21oi_1 _09326_ (.A1(_03235_),
    .A2(_02950_),
    .B1(_03236_),
    .Y(_03237_));
 sky130_fd_sc_hd__nand2_1 _09327_ (.A(_02785_),
    .B(_02821_),
    .Y(_03238_));
 sky130_fd_sc_hd__nand2_1 _09328_ (.A(_02905_),
    .B(_03238_),
    .Y(_03239_));
 sky130_fd_sc_hd__a21oi_1 _09329_ (.A1(_02783_),
    .A2(_02213_),
    .B1(_02897_),
    .Y(_03240_));
 sky130_fd_sc_hd__nand2_1 _09330_ (.A(_02687_),
    .B(_02895_),
    .Y(_03241_));
 sky130_fd_sc_hd__nand2_1 _09331_ (.A(_03240_),
    .B(_03241_),
    .Y(_03242_));
 sky130_fd_sc_hd__nand2_1 _09332_ (.A(_02963_),
    .B(_02734_),
    .Y(_03243_));
 sky130_fd_sc_hd__nand3_1 _09333_ (.A(_03239_),
    .B(_03242_),
    .C(_03243_),
    .Y(_03244_));
 sky130_fd_sc_hd__a21oi_1 _09334_ (.A1(_02783_),
    .A2(_02213_),
    .B1(_02904_),
    .Y(_03245_));
 sky130_fd_sc_hd__nand2_1 _09335_ (.A(_02898_),
    .B(_03245_),
    .Y(_03246_));
 sky130_fd_sc_hd__inv_2 _09336_ (.A(_03243_),
    .Y(_03247_));
 sky130_fd_sc_hd__nand2_1 _09337_ (.A(_03241_),
    .B(_03238_),
    .Y(_03248_));
 sky130_fd_sc_hd__nand3_1 _09338_ (.A(_03246_),
    .B(_03247_),
    .C(_03248_),
    .Y(_03249_));
 sky130_fd_sc_hd__nand2_1 _09339_ (.A(_03244_),
    .B(_03249_),
    .Y(_03250_));
 sky130_fd_sc_hd__nor2_1 _09340_ (.A(_02823_),
    .B(_03241_),
    .Y(_03251_));
 sky130_fd_sc_hd__a21oi_2 _09341_ (.A1(_02908_),
    .A2(_02907_),
    .B1(_03251_),
    .Y(_03252_));
 sky130_fd_sc_hd__inv_2 _09342_ (.A(_03252_),
    .Y(_03253_));
 sky130_fd_sc_hd__nand2_1 _09343_ (.A(_03250_),
    .B(_03253_),
    .Y(_03254_));
 sky130_fd_sc_hd__nand3_1 _09344_ (.A(_03252_),
    .B(_03244_),
    .C(_03249_),
    .Y(_03255_));
 sky130_fd_sc_hd__nand2_1 _09345_ (.A(_03254_),
    .B(_03255_),
    .Y(_03256_));
 sky130_fd_sc_hd__nor2_1 _09346_ (.A(_03051_),
    .B(_02578_),
    .Y(_03257_));
 sky130_fd_sc_hd__inv_2 _09347_ (.A(_03257_),
    .Y(_03258_));
 sky130_fd_sc_hd__nor2_1 _09348_ (.A(_03205_),
    .B(_03258_),
    .Y(_03259_));
 sky130_fd_sc_hd__nand2_1 _09349_ (.A(_03256_),
    .B(_03259_),
    .Y(_03260_));
 sky130_fd_sc_hd__inv_2 _09350_ (.A(_03259_),
    .Y(_03261_));
 sky130_fd_sc_hd__nand3_1 _09351_ (.A(_03254_),
    .B(_03255_),
    .C(_03261_),
    .Y(_03262_));
 sky130_fd_sc_hd__nand2_1 _09352_ (.A(_03260_),
    .B(_03262_),
    .Y(_03263_));
 sky130_fd_sc_hd__nor2_1 _09353_ (.A(_03237_),
    .B(_03263_),
    .Y(_03264_));
 sky130_fd_sc_hd__nand2_1 _09354_ (.A(_03263_),
    .B(_03237_),
    .Y(_03265_));
 sky130_fd_sc_hd__nand2b_1 _09355_ (.A_N(_03264_),
    .B(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__nand2_1 _09356_ (.A(_03266_),
    .B(_02954_),
    .Y(_03267_));
 sky130_fd_sc_hd__inv_2 _09357_ (.A(_03265_),
    .Y(_03268_));
 sky130_fd_sc_hd__nor2_1 _09358_ (.A(_03264_),
    .B(_03268_),
    .Y(_03269_));
 sky130_fd_sc_hd__nor2_1 _09359_ (.A(_02828_),
    .B(_02955_),
    .Y(_03270_));
 sky130_fd_sc_hd__nand2_1 _09360_ (.A(_03269_),
    .B(_03270_),
    .Y(_03271_));
 sky130_fd_sc_hd__inv_2 _09361_ (.A(_03224_),
    .Y(_03272_));
 sky130_fd_sc_hd__a21o_1 _09362_ (.A1(_03267_),
    .A2(_03271_),
    .B1(_03272_),
    .X(_03273_));
 sky130_fd_sc_hd__clkbuf_4 _09363_ (.A(_03079_),
    .X(_03274_));
 sky130_fd_sc_hd__nand3_1 _09364_ (.A(_03267_),
    .B(_03272_),
    .C(_03271_),
    .Y(_03275_));
 sky130_fd_sc_hd__nand3_1 _09365_ (.A(_03273_),
    .B(_03274_),
    .C(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__nand3_1 _09366_ (.A(_03234_),
    .B(_03276_),
    .C(_00622_),
    .Y(_03277_));
 sky130_fd_sc_hd__nand2_1 _09367_ (.A(_03206_),
    .B(_00549_),
    .Y(_03278_));
 sky130_fd_sc_hd__nand2_1 _09368_ (.A(_03277_),
    .B(_03278_),
    .Y(_03279_));
 sky130_fd_sc_hd__and3_1 _09369_ (.A(_00620_),
    .B(_00523_),
    .C(_00582_),
    .X(_03280_));
 sky130_fd_sc_hd__nand2_1 _09370_ (.A(_03280_),
    .B(\Add.sub ),
    .Y(_03281_));
 sky130_fd_sc_hd__nand2_1 _09371_ (.A(_03279_),
    .B(_03281_),
    .Y(_03282_));
 sky130_fd_sc_hd__inv_2 _09372_ (.A(_03281_),
    .Y(_03283_));
 sky130_fd_sc_hd__nand3_1 _09373_ (.A(_03277_),
    .B(_03278_),
    .C(_03283_),
    .Y(_03284_));
 sky130_fd_sc_hd__nand2_1 _09374_ (.A(_03282_),
    .B(_03284_),
    .Y(_03285_));
 sky130_fd_sc_hd__a21oi_1 _09375_ (.A1(_02985_),
    .A2(_02982_),
    .B1(_03233_),
    .Y(_03286_));
 sky130_fd_sc_hd__inv_2 _09376_ (.A(_03286_),
    .Y(_03287_));
 sky130_fd_sc_hd__nand2_1 _09377_ (.A(_03285_),
    .B(_03287_),
    .Y(_03288_));
 sky130_fd_sc_hd__nand3_1 _09378_ (.A(_03286_),
    .B(_03282_),
    .C(_03284_),
    .Y(_03289_));
 sky130_fd_sc_hd__nand2_1 _09379_ (.A(_03288_),
    .B(_03289_),
    .Y(_03290_));
 sky130_fd_sc_hd__nor2_4 _09380_ (.A(_03046_),
    .B(_03290_),
    .Y(_03291_));
 sky130_fd_sc_hd__and2_1 _09381_ (.A(_03290_),
    .B(_03046_),
    .X(_03292_));
 sky130_fd_sc_hd__nor2_2 _09382_ (.A(_03291_),
    .B(_03292_),
    .Y(_03293_));
 sky130_fd_sc_hd__nor2_1 _09383_ (.A(_02653_),
    .B(_03293_),
    .Y(_03294_));
 sky130_fd_sc_hd__a211o_1 _09384_ (.A1(_00789_),
    .A2(_02654_),
    .B1(_02753_),
    .C1(_03294_),
    .X(_03295_));
 sky130_fd_sc_hd__inv_2 _09385_ (.A(_03295_),
    .Y(_00248_));
 sky130_fd_sc_hd__nor2_1 _09386_ (.A(_00536_),
    .B(_03280_),
    .Y(_03296_));
 sky130_fd_sc_hd__nand2_1 _09387_ (.A(_03279_),
    .B(_03296_),
    .Y(_03297_));
 sky130_fd_sc_hd__nand2_1 _09388_ (.A(_03289_),
    .B(_03297_),
    .Y(_03298_));
 sky130_fd_sc_hd__inv_2 _09389_ (.A(_03298_),
    .Y(_03299_));
 sky130_fd_sc_hd__o21bai_1 _09390_ (.A1(_02954_),
    .A2(_03268_),
    .B1_N(_03264_),
    .Y(_03300_));
 sky130_fd_sc_hd__a21oi_1 _09391_ (.A1(_02947_),
    .A2(_02237_),
    .B1(_02904_),
    .Y(_03301_));
 sky130_fd_sc_hd__nand2_1 _09392_ (.A(_03301_),
    .B(_03240_),
    .Y(_03302_));
 sky130_fd_sc_hd__nand2_1 _09393_ (.A(_02734_),
    .B(_03079_),
    .Y(_03303_));
 sky130_fd_sc_hd__inv_2 _09394_ (.A(_03303_),
    .Y(_03304_));
 sky130_fd_sc_hd__nand2_1 _09395_ (.A(_03304_),
    .B(_03019_),
    .Y(_03305_));
 sky130_fd_sc_hd__inv_2 _09396_ (.A(_03305_),
    .Y(_03306_));
 sky130_fd_sc_hd__nand2_1 _09397_ (.A(_02963_),
    .B(_02821_),
    .Y(_03307_));
 sky130_fd_sc_hd__nand2_1 _09398_ (.A(_02785_),
    .B(_02895_),
    .Y(_03308_));
 sky130_fd_sc_hd__nand2_1 _09399_ (.A(_03307_),
    .B(_03308_),
    .Y(_03309_));
 sky130_fd_sc_hd__nand3_1 _09400_ (.A(_03302_),
    .B(_03306_),
    .C(_03309_),
    .Y(_03310_));
 sky130_fd_sc_hd__nand3_1 _09401_ (.A(_03308_),
    .B(_02821_),
    .C(_02963_),
    .Y(_03311_));
 sky130_fd_sc_hd__nand2_1 _09402_ (.A(_03245_),
    .B(_03307_),
    .Y(_03312_));
 sky130_fd_sc_hd__nand3_1 _09403_ (.A(_03311_),
    .B(_03312_),
    .C(_03305_),
    .Y(_03313_));
 sky130_fd_sc_hd__nand2_1 _09404_ (.A(_03310_),
    .B(_03313_),
    .Y(_03314_));
 sky130_fd_sc_hd__nor2_1 _09405_ (.A(_02822_),
    .B(_03308_),
    .Y(_03315_));
 sky130_fd_sc_hd__a21oi_2 _09406_ (.A1(_03248_),
    .A2(_03247_),
    .B1(_03315_),
    .Y(_03316_));
 sky130_fd_sc_hd__inv_2 _09407_ (.A(_03316_),
    .Y(_03317_));
 sky130_fd_sc_hd__nand2_1 _09408_ (.A(_03314_),
    .B(_03317_),
    .Y(_03318_));
 sky130_fd_sc_hd__nand3_1 _09409_ (.A(_03316_),
    .B(_03310_),
    .C(_03313_),
    .Y(_03319_));
 sky130_fd_sc_hd__nand2_1 _09410_ (.A(_03318_),
    .B(_03319_),
    .Y(_03320_));
 sky130_fd_sc_hd__nand2_1 _09411_ (.A(_02611_),
    .B(\Qset[1][5] ),
    .Y(_03321_));
 sky130_fd_sc_hd__nand2_1 _09412_ (.A(_03321_),
    .B(_02591_),
    .Y(_03322_));
 sky130_fd_sc_hd__nand2_1 _09413_ (.A(_02582_),
    .B(\Qset[0][5] ),
    .Y(_03323_));
 sky130_fd_sc_hd__inv_2 _09414_ (.A(_03323_),
    .Y(_03324_));
 sky130_fd_sc_hd__nand2_1 _09415_ (.A(_02582_),
    .B(\Qset[2][5] ),
    .Y(_03325_));
 sky130_fd_sc_hd__nand2_1 _09416_ (.A(_02992_),
    .B(\Qset[3][5] ),
    .Y(_03326_));
 sky130_fd_sc_hd__nand3_1 _09417_ (.A(_03325_),
    .B(_02991_),
    .C(_03326_),
    .Y(_03327_));
 sky130_fd_sc_hd__o21ai_2 _09418_ (.A1(_03322_),
    .A2(_03324_),
    .B1(_03327_),
    .Y(_03328_));
 sky130_fd_sc_hd__nand2_1 _09419_ (.A(_03328_),
    .B(_00581_),
    .Y(_03329_));
 sky130_fd_sc_hd__nand2_1 _09420_ (.A(_02273_),
    .B(_02161_),
    .Y(_03330_));
 sky130_fd_sc_hd__nand3_1 _09421_ (.A(_03329_),
    .B(_03330_),
    .C(_02540_),
    .Y(_03331_));
 sky130_fd_sc_hd__nand2_1 _09422_ (.A(_03001_),
    .B(\Oset[3][5] ),
    .Y(_03332_));
 sky130_fd_sc_hd__o211ai_2 _09423_ (.A1(_03001_),
    .A2(_02274_),
    .B1(_02991_),
    .C1(_03332_),
    .Y(_03333_));
 sky130_fd_sc_hd__nand2_1 _09424_ (.A(_03001_),
    .B(\Oset[1][5] ),
    .Y(_03334_));
 sky130_fd_sc_hd__o211ai_2 _09425_ (.A1(_02992_),
    .A2(_02277_),
    .B1(_03004_),
    .C1(_03334_),
    .Y(_03335_));
 sky130_fd_sc_hd__nand3_1 _09426_ (.A(_03333_),
    .B(_03335_),
    .C(_02551_),
    .Y(_03336_));
 sky130_fd_sc_hd__nand3_1 _09427_ (.A(_03331_),
    .B(_01155_),
    .C(_03336_),
    .Y(_03337_));
 sky130_fd_sc_hd__nand2_1 _09428_ (.A(_02280_),
    .B(_00583_),
    .Y(_03338_));
 sky130_fd_sc_hd__nand2_1 _09429_ (.A(_03337_),
    .B(_03338_),
    .Y(_03339_));
 sky130_fd_sc_hd__nand2_1 _09430_ (.A(_03339_),
    .B(_02556_),
    .Y(_03340_));
 sky130_fd_sc_hd__buf_6 _09431_ (.A(_02582_),
    .X(_03341_));
 sky130_fd_sc_hd__nand2_1 _09432_ (.A(_03341_),
    .B(_02281_),
    .Y(_03342_));
 sky130_fd_sc_hd__o21a_1 _09433_ (.A1(\H[1][5] ),
    .A2(_03341_),
    .B1(_02591_),
    .X(_03343_));
 sky130_fd_sc_hd__mux2_1 _09434_ (.A0(\H[2][5] ),
    .A1(\H[3][5] ),
    .S(_02611_),
    .X(_03344_));
 sky130_fd_sc_hd__buf_4 _09435_ (.A(_02991_),
    .X(_03345_));
 sky130_fd_sc_hd__a22oi_4 _09436_ (.A1(_03342_),
    .A2(_03343_),
    .B1(_03344_),
    .B2(_03345_),
    .Y(_03346_));
 sky130_fd_sc_hd__a21oi_1 _09437_ (.A1(_03346_),
    .A2(_02572_),
    .B1(_00587_),
    .Y(_03347_));
 sky130_fd_sc_hd__nand2_2 _09438_ (.A(_03340_),
    .B(_03347_),
    .Y(_03348_));
 sky130_fd_sc_hd__nand2_2 _09439_ (.A(_03348_),
    .B(_02286_),
    .Y(_03349_));
 sky130_fd_sc_hd__inv_2 _09440_ (.A(_03349_),
    .Y(_03350_));
 sky130_fd_sc_hd__nor2_1 _09441_ (.A(_03350_),
    .B(_03258_),
    .Y(_03351_));
 sky130_fd_sc_hd__nand2_1 _09442_ (.A(_03320_),
    .B(_03351_),
    .Y(_03352_));
 sky130_fd_sc_hd__nand3b_1 _09443_ (.A_N(_03351_),
    .B(_03318_),
    .C(_03319_),
    .Y(_03353_));
 sky130_fd_sc_hd__nand2_1 _09444_ (.A(_03352_),
    .B(_03353_),
    .Y(_03354_));
 sky130_fd_sc_hd__nand2_1 _09445_ (.A(_03250_),
    .B(_03252_),
    .Y(_03355_));
 sky130_fd_sc_hd__nor2_1 _09446_ (.A(_03252_),
    .B(_03250_),
    .Y(_03356_));
 sky130_fd_sc_hd__a21oi_2 _09447_ (.A1(_03355_),
    .A2(_03259_),
    .B1(_03356_),
    .Y(_03357_));
 sky130_fd_sc_hd__inv_2 _09448_ (.A(_03357_),
    .Y(_03358_));
 sky130_fd_sc_hd__nand2_1 _09449_ (.A(_03354_),
    .B(_03358_),
    .Y(_03359_));
 sky130_fd_sc_hd__nand3_1 _09450_ (.A(_03357_),
    .B(_03352_),
    .C(_03353_),
    .Y(_03360_));
 sky130_fd_sc_hd__nand2_1 _09451_ (.A(_03359_),
    .B(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hd__nand2_1 _09452_ (.A(_03300_),
    .B(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__a21oi_1 _09453_ (.A1(_03270_),
    .A2(_03265_),
    .B1(_03264_),
    .Y(_03363_));
 sky130_fd_sc_hd__inv_2 _09454_ (.A(_03361_),
    .Y(_03364_));
 sky130_fd_sc_hd__nand2_1 _09455_ (.A(_03363_),
    .B(_03364_),
    .Y(_03365_));
 sky130_fd_sc_hd__nand2_1 _09456_ (.A(_03362_),
    .B(_03365_),
    .Y(_03366_));
 sky130_fd_sc_hd__a21bo_1 _09457_ (.A1(_03176_),
    .A2(_03052_),
    .B1_N(_03220_),
    .X(_03367_));
 sky130_fd_sc_hd__inv_2 _09458_ (.A(_03367_),
    .Y(_03368_));
 sky130_fd_sc_hd__nor2_1 _09459_ (.A(_03225_),
    .B(_03368_),
    .Y(_03369_));
 sky130_fd_sc_hd__nand2_1 _09460_ (.A(_03366_),
    .B(_03369_),
    .Y(_03370_));
 sky130_fd_sc_hd__inv_2 _09461_ (.A(_03369_),
    .Y(_03371_));
 sky130_fd_sc_hd__nand3_1 _09462_ (.A(_03362_),
    .B(_03365_),
    .C(_03371_),
    .Y(_03372_));
 sky130_fd_sc_hd__nand3_1 _09463_ (.A(_03370_),
    .B(_03275_),
    .C(_03372_),
    .Y(_03373_));
 sky130_fd_sc_hd__nand2_1 _09464_ (.A(_03366_),
    .B(_03371_),
    .Y(_03374_));
 sky130_fd_sc_hd__inv_2 _09465_ (.A(_03275_),
    .Y(_03375_));
 sky130_fd_sc_hd__nand3_1 _09466_ (.A(_03362_),
    .B(_03365_),
    .C(_03369_),
    .Y(_03376_));
 sky130_fd_sc_hd__nand3_1 _09467_ (.A(_03374_),
    .B(_03375_),
    .C(_03376_),
    .Y(_03377_));
 sky130_fd_sc_hd__nand2_1 _09468_ (.A(_03373_),
    .B(_03377_),
    .Y(_03378_));
 sky130_fd_sc_hd__nand2_1 _09469_ (.A(_03378_),
    .B(_03274_),
    .Y(_03379_));
 sky130_fd_sc_hd__o21bai_1 _09470_ (.A1(_03228_),
    .A2(_03216_),
    .B1_N(_03214_),
    .Y(_03380_));
 sky130_fd_sc_hd__a21boi_2 _09471_ (.A1(_03207_),
    .A2(_03211_),
    .B1_N(_03210_),
    .Y(_03381_));
 sky130_fd_sc_hd__inv_2 _09472_ (.A(_03381_),
    .Y(_03382_));
 sky130_fd_sc_hd__inv_2 _09473_ (.A(_03145_),
    .Y(_03383_));
 sky130_fd_sc_hd__nor2_1 _09474_ (.A(_03205_),
    .B(_03383_),
    .Y(_03384_));
 sky130_fd_sc_hd__nand2_1 _09475_ (.A(_03184_),
    .B(_03076_),
    .Y(_03385_));
 sky130_fd_sc_hd__nor2_1 _09476_ (.A(_03190_),
    .B(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__nand2_1 _09477_ (.A(_03184_),
    .B(_03110_),
    .Y(_03387_));
 sky130_fd_sc_hd__nand2_1 _09478_ (.A(_03116_),
    .B(_03076_),
    .Y(_03388_));
 sky130_fd_sc_hd__nand2_1 _09479_ (.A(_03387_),
    .B(_03388_),
    .Y(_03389_));
 sky130_fd_sc_hd__inv_2 _09480_ (.A(_03389_),
    .Y(_03390_));
 sky130_fd_sc_hd__nor2_1 _09481_ (.A(_03386_),
    .B(_03390_),
    .Y(_03391_));
 sky130_fd_sc_hd__or2_1 _09482_ (.A(_03384_),
    .B(_03391_),
    .X(_03392_));
 sky130_fd_sc_hd__nand2_1 _09483_ (.A(_03391_),
    .B(_03384_),
    .Y(_03393_));
 sky130_fd_sc_hd__nand2_1 _09484_ (.A(_03392_),
    .B(_03393_),
    .Y(_03394_));
 sky130_fd_sc_hd__a21oi_2 _09485_ (.A1(_03192_),
    .A2(_03197_),
    .B1(_03191_),
    .Y(_03395_));
 sky130_fd_sc_hd__inv_2 _09486_ (.A(_03395_),
    .Y(_03396_));
 sky130_fd_sc_hd__nand2_1 _09487_ (.A(_03394_),
    .B(_03396_),
    .Y(_03397_));
 sky130_fd_sc_hd__nand3_1 _09488_ (.A(_03392_),
    .B(_03395_),
    .C(_03393_),
    .Y(_03398_));
 sky130_fd_sc_hd__nand2_1 _09489_ (.A(_03397_),
    .B(_03398_),
    .Y(_03399_));
 sky130_fd_sc_hd__nor2_1 _09490_ (.A(_03350_),
    .B(_03206_),
    .Y(_03400_));
 sky130_fd_sc_hd__nand2_1 _09491_ (.A(_03399_),
    .B(_03400_),
    .Y(_03401_));
 sky130_fd_sc_hd__nand3b_1 _09492_ (.A_N(_03400_),
    .B(_03397_),
    .C(_03398_),
    .Y(_03402_));
 sky130_fd_sc_hd__nand2_1 _09493_ (.A(_03401_),
    .B(_03402_),
    .Y(_03403_));
 sky130_fd_sc_hd__nand2_1 _09494_ (.A(_03382_),
    .B(_03403_),
    .Y(_03404_));
 sky130_fd_sc_hd__nand3_1 _09495_ (.A(_03381_),
    .B(_03402_),
    .C(_03401_),
    .Y(_03405_));
 sky130_fd_sc_hd__nand2_1 _09496_ (.A(_03404_),
    .B(_03405_),
    .Y(_03406_));
 sky130_fd_sc_hd__nand2_1 _09497_ (.A(_03380_),
    .B(_03406_),
    .Y(_03407_));
 sky130_fd_sc_hd__a21oi_1 _09498_ (.A1(_03231_),
    .A2(_03215_),
    .B1(_03214_),
    .Y(_03408_));
 sky130_fd_sc_hd__inv_2 _09499_ (.A(_03406_),
    .Y(_03409_));
 sky130_fd_sc_hd__nand2_1 _09500_ (.A(_03408_),
    .B(_03409_),
    .Y(_03410_));
 sky130_fd_sc_hd__nand2_2 _09501_ (.A(_03407_),
    .B(_03410_),
    .Y(_03411_));
 sky130_fd_sc_hd__nand2_1 _09502_ (.A(_03411_),
    .B(_03233_),
    .Y(_03412_));
 sky130_fd_sc_hd__nand3_1 _09503_ (.A(_03379_),
    .B(_00623_),
    .C(_03412_),
    .Y(_03413_));
 sky130_fd_sc_hd__nand2_1 _09504_ (.A(_03145_),
    .B(_00556_),
    .Y(_03414_));
 sky130_fd_sc_hd__nand3_1 _09505_ (.A(_03413_),
    .B(_02092_),
    .C(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__nand3_1 _09506_ (.A(_03373_),
    .B(_03377_),
    .C(_03274_),
    .Y(_03416_));
 sky130_fd_sc_hd__nand3_1 _09507_ (.A(_03407_),
    .B(_03410_),
    .C(_03233_),
    .Y(_03417_));
 sky130_fd_sc_hd__nand3_1 _09508_ (.A(_03416_),
    .B(_00623_),
    .C(_03417_),
    .Y(_03418_));
 sky130_fd_sc_hd__nand2_1 _09509_ (.A(_03383_),
    .B(_00556_),
    .Y(_03419_));
 sky130_fd_sc_hd__nand3_1 _09510_ (.A(_03418_),
    .B(_00536_),
    .C(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__buf_6 _09511_ (.A(_03349_),
    .X(_03421_));
 sky130_fd_sc_hd__a21o_1 _09512_ (.A1(\H[3][5] ),
    .A2(_03033_),
    .B1(_03026_),
    .X(_03422_));
 sky130_fd_sc_hd__a21o_1 _09513_ (.A1(\H[2][5] ),
    .A2(_03022_),
    .B1(_03422_),
    .X(_03423_));
 sky130_fd_sc_hd__nor2_1 _09514_ (.A(_03033_),
    .B(_02281_),
    .Y(_03424_));
 sky130_fd_sc_hd__a211o_1 _09515_ (.A1(\H[1][5] ),
    .A2(_03033_),
    .B1(_02840_),
    .C1(_03424_),
    .X(_03425_));
 sky130_fd_sc_hd__nand2_1 _09516_ (.A(_03021_),
    .B(\Oset[0][5] ),
    .Y(_03426_));
 sky130_fd_sc_hd__nand2_1 _09517_ (.A(\Oset[1][5] ),
    .B(_03024_),
    .Y(_03427_));
 sky130_fd_sc_hd__a21oi_1 _09518_ (.A1(\Oset[3][5] ),
    .A2(_03024_),
    .B1(_02837_),
    .Y(_03428_));
 sky130_fd_sc_hd__nand2_1 _09519_ (.A(_03021_),
    .B(\Oset[2][5] ),
    .Y(_03429_));
 sky130_fd_sc_hd__a32o_1 _09520_ (.A1(_03426_),
    .A2(_03427_),
    .A3(_03026_),
    .B1(_03428_),
    .B2(_03429_),
    .X(_03430_));
 sky130_fd_sc_hd__nand2_1 _09521_ (.A(_02632_),
    .B(\Qset[0][5] ),
    .Y(_03431_));
 sky130_fd_sc_hd__nand2_1 _09522_ (.A(\Qset[1][5] ),
    .B(_03024_),
    .Y(_03432_));
 sky130_fd_sc_hd__a21oi_1 _09523_ (.A1(\Qset[3][5] ),
    .A2(_03024_),
    .B1(_02837_),
    .Y(_03433_));
 sky130_fd_sc_hd__nand2_1 _09524_ (.A(_03021_),
    .B(\Qset[2][5] ),
    .Y(_03434_));
 sky130_fd_sc_hd__a32o_1 _09525_ (.A1(_03431_),
    .A2(_03432_),
    .A3(_02837_),
    .B1(_03433_),
    .B2(_03434_),
    .X(_03435_));
 sky130_fd_sc_hd__mux2_1 _09526_ (.A0(_03430_),
    .A1(_03435_),
    .S(_00646_),
    .X(_03436_));
 sky130_fd_sc_hd__nor2_1 _09527_ (.A(_01536_),
    .B(_03436_),
    .Y(_03437_));
 sky130_fd_sc_hd__a311o_2 _09528_ (.A1(_01536_),
    .A2(_03423_),
    .A3(_03425_),
    .B1(_00549_),
    .C1(_03437_),
    .X(_03438_));
 sky130_fd_sc_hd__o21ai_2 _09529_ (.A1(_00623_),
    .A2(_03421_),
    .B1(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__nand3_1 _09530_ (.A(_03415_),
    .B(_03420_),
    .C(_03439_),
    .Y(_03440_));
 sky130_fd_sc_hd__nand3_1 _09531_ (.A(_03413_),
    .B(_00536_),
    .C(_03414_),
    .Y(_03441_));
 sky130_fd_sc_hd__nand3_1 _09532_ (.A(_03418_),
    .B(_02092_),
    .C(_03419_),
    .Y(_03442_));
 sky130_fd_sc_hd__inv_2 _09533_ (.A(_03439_),
    .Y(_03443_));
 sky130_fd_sc_hd__nand3_1 _09534_ (.A(_03441_),
    .B(_03442_),
    .C(_03443_),
    .Y(_03444_));
 sky130_fd_sc_hd__nand2_1 _09535_ (.A(_03440_),
    .B(_03444_),
    .Y(_03445_));
 sky130_fd_sc_hd__nor2_1 _09536_ (.A(_03299_),
    .B(_03445_),
    .Y(_03446_));
 sky130_fd_sc_hd__nand2_1 _09537_ (.A(_03445_),
    .B(_03299_),
    .Y(_03447_));
 sky130_fd_sc_hd__or2b_2 _09538_ (.A(_03446_),
    .B_N(_03447_),
    .X(_03448_));
 sky130_fd_sc_hd__xnor2_4 _09539_ (.A(_03291_),
    .B(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__nor2_1 _09540_ (.A(_02653_),
    .B(_03449_),
    .Y(_03450_));
 sky130_fd_sc_hd__a211o_1 _09541_ (.A1(_00812_),
    .A2(_02654_),
    .B1(_02753_),
    .C1(_03450_),
    .X(_03451_));
 sky130_fd_sc_hd__inv_2 _09542_ (.A(_03451_),
    .Y(_00249_));
 sky130_fd_sc_hd__a21oi_4 _09543_ (.A1(_03447_),
    .A2(_03291_),
    .B1(_03446_),
    .Y(_03452_));
 sky130_fd_sc_hd__nand3_1 _09544_ (.A(_03269_),
    .B(_03270_),
    .C(_03361_),
    .Y(_03453_));
 sky130_fd_sc_hd__nand2_1 _09545_ (.A(_03354_),
    .B(_03357_),
    .Y(_03454_));
 sky130_fd_sc_hd__nor2_1 _09546_ (.A(_03357_),
    .B(_03354_),
    .Y(_03455_));
 sky130_fd_sc_hd__a21oi_1 _09547_ (.A1(_03264_),
    .A2(_03454_),
    .B1(_03455_),
    .Y(_03456_));
 sky130_fd_sc_hd__nand2_1 _09548_ (.A(_03453_),
    .B(_03456_),
    .Y(_03457_));
 sky130_fd_sc_hd__nand2_1 _09549_ (.A(_02821_),
    .B(_03079_),
    .Y(_03458_));
 sky130_fd_sc_hd__a21oi_1 _09550_ (.A1(_03018_),
    .A2(_02264_),
    .B1(_03458_),
    .Y(_03459_));
 sky130_fd_sc_hd__nand2_1 _09551_ (.A(_03459_),
    .B(_03301_),
    .Y(_03460_));
 sky130_fd_sc_hd__a21oi_1 _09552_ (.A1(_03348_),
    .A2(_02286_),
    .B1(_03303_),
    .Y(_03461_));
 sky130_fd_sc_hd__inv_2 _09553_ (.A(_03458_),
    .Y(_03462_));
 sky130_fd_sc_hd__nand2_1 _09554_ (.A(_03020_),
    .B(_03462_),
    .Y(_03463_));
 sky130_fd_sc_hd__nand2_1 _09555_ (.A(_02963_),
    .B(_02895_),
    .Y(_03464_));
 sky130_fd_sc_hd__nand2_1 _09556_ (.A(_03463_),
    .B(_03464_),
    .Y(_03465_));
 sky130_fd_sc_hd__nand3_1 _09557_ (.A(_03460_),
    .B(_03461_),
    .C(_03465_),
    .Y(_03466_));
 sky130_fd_sc_hd__nand2_1 _09558_ (.A(_03459_),
    .B(_03464_),
    .Y(_03467_));
 sky130_fd_sc_hd__nand2_1 _09559_ (.A(_03463_),
    .B(_03301_),
    .Y(_03468_));
 sky130_fd_sc_hd__nand2_1 _09560_ (.A(_03421_),
    .B(_03304_),
    .Y(_03469_));
 sky130_fd_sc_hd__nand3_1 _09561_ (.A(_03467_),
    .B(_03468_),
    .C(_03469_),
    .Y(_03470_));
 sky130_fd_sc_hd__nand2_1 _09562_ (.A(_03466_),
    .B(_03470_),
    .Y(_03471_));
 sky130_fd_sc_hd__nor2_1 _09563_ (.A(_03238_),
    .B(_03464_),
    .Y(_03472_));
 sky130_fd_sc_hd__a21oi_2 _09564_ (.A1(_03306_),
    .A2(_03309_),
    .B1(_03472_),
    .Y(_03473_));
 sky130_fd_sc_hd__inv_2 _09565_ (.A(_03473_),
    .Y(_03474_));
 sky130_fd_sc_hd__nand2_1 _09566_ (.A(_03471_),
    .B(_03474_),
    .Y(_03475_));
 sky130_fd_sc_hd__nand3_1 _09567_ (.A(_03473_),
    .B(_03466_),
    .C(_03470_),
    .Y(_03476_));
 sky130_fd_sc_hd__nand2_1 _09568_ (.A(_03475_),
    .B(_03476_),
    .Y(_03477_));
 sky130_fd_sc_hd__nor2_1 _09569_ (.A(_02611_),
    .B(_02299_),
    .Y(_03478_));
 sky130_fd_sc_hd__a21o_1 _09570_ (.A1(_02586_),
    .A2(\Oset[1][6] ),
    .B1(_02584_),
    .X(_03479_));
 sky130_fd_sc_hd__nand2_1 _09571_ (.A(_02611_),
    .B(\Oset[3][6] ),
    .Y(_03480_));
 sky130_fd_sc_hd__o211ai_1 _09572_ (.A1(_02611_),
    .A2(_02296_),
    .B1(_02584_),
    .C1(_03480_),
    .Y(_03481_));
 sky130_fd_sc_hd__o21ai_2 _09573_ (.A1(_03478_),
    .A2(_03479_),
    .B1(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__o21ai_1 _09574_ (.A1(_02540_),
    .A2(_03482_),
    .B1(_01154_),
    .Y(_03483_));
 sky130_fd_sc_hd__inv_2 _09575_ (.A(_03483_),
    .Y(_03484_));
 sky130_fd_sc_hd__nor2_1 _09576_ (.A(_02992_),
    .B(_02292_),
    .Y(_03485_));
 sky130_fd_sc_hd__a21o_1 _09577_ (.A1(_02992_),
    .A2(\Qset[1][6] ),
    .B1(_02991_),
    .X(_03486_));
 sky130_fd_sc_hd__nand2_1 _09578_ (.A(_03001_),
    .B(\Qset[3][6] ),
    .Y(_03487_));
 sky130_fd_sc_hd__o211ai_1 _09579_ (.A1(_03001_),
    .A2(_02289_),
    .B1(_02991_),
    .C1(_03487_),
    .Y(_03488_));
 sky130_fd_sc_hd__o21ai_2 _09580_ (.A1(_03485_),
    .A2(_03486_),
    .B1(_03488_),
    .Y(_03489_));
 sky130_fd_sc_hd__nand2_1 _09581_ (.A(_03489_),
    .B(_00581_),
    .Y(_03490_));
 sky130_fd_sc_hd__nand2_1 _09582_ (.A(_02295_),
    .B(_02161_),
    .Y(_03491_));
 sky130_fd_sc_hd__nand3_1 _09583_ (.A(_03490_),
    .B(_03491_),
    .C(_02540_),
    .Y(_03492_));
 sky130_fd_sc_hd__nand2_1 _09584_ (.A(_03484_),
    .B(_03492_),
    .Y(_03493_));
 sky130_fd_sc_hd__nand2_1 _09585_ (.A(_02302_),
    .B(_00584_),
    .Y(_03494_));
 sky130_fd_sc_hd__nand2_1 _09586_ (.A(_03493_),
    .B(_03494_),
    .Y(_03495_));
 sky130_fd_sc_hd__nand2_1 _09587_ (.A(_03495_),
    .B(_02556_),
    .Y(_03496_));
 sky130_fd_sc_hd__nand2_1 _09588_ (.A(_03341_),
    .B(\H[2][6] ),
    .Y(_03497_));
 sky130_fd_sc_hd__buf_6 _09589_ (.A(_02992_),
    .X(_03498_));
 sky130_fd_sc_hd__nand2_1 _09590_ (.A(_03498_),
    .B(\H[3][6] ),
    .Y(_03499_));
 sky130_fd_sc_hd__nand2_1 _09591_ (.A(_03001_),
    .B(\H[1][6] ),
    .Y(_03500_));
 sky130_fd_sc_hd__o211a_1 _09592_ (.A1(_02992_),
    .A2(_02303_),
    .B1(_03004_),
    .C1(_03500_),
    .X(_03501_));
 sky130_fd_sc_hd__a31o_2 _09593_ (.A1(_03345_),
    .A2(_03497_),
    .A3(_03499_),
    .B1(_03501_),
    .X(_03502_));
 sky130_fd_sc_hd__a21oi_1 _09594_ (.A1(_03502_),
    .A2(_02573_),
    .B1(_00587_),
    .Y(_03503_));
 sky130_fd_sc_hd__nand2_2 _09595_ (.A(_03496_),
    .B(_03503_),
    .Y(_03504_));
 sky130_fd_sc_hd__nand2_2 _09596_ (.A(_03504_),
    .B(_02308_),
    .Y(_03505_));
 sky130_fd_sc_hd__buf_6 _09597_ (.A(_03505_),
    .X(_03506_));
 sky130_fd_sc_hd__inv_2 _09598_ (.A(_03506_),
    .Y(_03507_));
 sky130_fd_sc_hd__nor2_1 _09599_ (.A(_03507_),
    .B(_03258_),
    .Y(_03508_));
 sky130_fd_sc_hd__nand2_1 _09600_ (.A(_03477_),
    .B(_03508_),
    .Y(_03509_));
 sky130_fd_sc_hd__nand3b_1 _09601_ (.A_N(_03508_),
    .B(_03475_),
    .C(_03476_),
    .Y(_03510_));
 sky130_fd_sc_hd__nand2_1 _09602_ (.A(_03509_),
    .B(_03510_),
    .Y(_03511_));
 sky130_fd_sc_hd__nand2_1 _09603_ (.A(_03314_),
    .B(_03316_),
    .Y(_03512_));
 sky130_fd_sc_hd__nor2_1 _09604_ (.A(_03316_),
    .B(_03314_),
    .Y(_03513_));
 sky130_fd_sc_hd__a21oi_2 _09605_ (.A1(_03512_),
    .A2(_03351_),
    .B1(_03513_),
    .Y(_03514_));
 sky130_fd_sc_hd__inv_2 _09606_ (.A(_03514_),
    .Y(_03515_));
 sky130_fd_sc_hd__nand2_1 _09607_ (.A(_03511_),
    .B(_03515_),
    .Y(_03516_));
 sky130_fd_sc_hd__nand3_1 _09608_ (.A(_03514_),
    .B(_03509_),
    .C(_03510_),
    .Y(_03517_));
 sky130_fd_sc_hd__nand2_1 _09609_ (.A(_03516_),
    .B(_03517_),
    .Y(_03518_));
 sky130_fd_sc_hd__nand2_1 _09610_ (.A(_03457_),
    .B(_03518_),
    .Y(_03519_));
 sky130_fd_sc_hd__nand3b_1 _09611_ (.A_N(_03518_),
    .B(_03453_),
    .C(_03456_),
    .Y(_03520_));
 sky130_fd_sc_hd__nand2_1 _09612_ (.A(_03519_),
    .B(_03520_),
    .Y(_03521_));
 sky130_fd_sc_hd__or2_1 _09613_ (.A(_03225_),
    .B(_03223_),
    .X(_03522_));
 sky130_fd_sc_hd__nand2_1 _09614_ (.A(_03522_),
    .B(_03226_),
    .Y(_03523_));
 sky130_fd_sc_hd__inv_2 _09615_ (.A(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__nand2_1 _09616_ (.A(_03521_),
    .B(_03524_),
    .Y(_03525_));
 sky130_fd_sc_hd__nand3_1 _09617_ (.A(_03519_),
    .B(_03520_),
    .C(_03523_),
    .Y(_03526_));
 sky130_fd_sc_hd__nand2_1 _09618_ (.A(_03525_),
    .B(_03526_),
    .Y(_03527_));
 sky130_fd_sc_hd__nand2_1 _09619_ (.A(_03377_),
    .B(_03376_),
    .Y(_03528_));
 sky130_fd_sc_hd__nand2_1 _09620_ (.A(_03527_),
    .B(_03528_),
    .Y(_03529_));
 sky130_fd_sc_hd__nand2_1 _09621_ (.A(_03521_),
    .B(_03523_),
    .Y(_03530_));
 sky130_fd_sc_hd__nand3_1 _09622_ (.A(_03519_),
    .B(_03520_),
    .C(_03524_),
    .Y(_03531_));
 sky130_fd_sc_hd__nand2_1 _09623_ (.A(_03530_),
    .B(_03531_),
    .Y(_03532_));
 sky130_fd_sc_hd__a21boi_1 _09624_ (.A1(_03374_),
    .A2(_03375_),
    .B1_N(_03376_),
    .Y(_03533_));
 sky130_fd_sc_hd__nand2_1 _09625_ (.A(_03532_),
    .B(_03533_),
    .Y(_03534_));
 sky130_fd_sc_hd__nand2_1 _09626_ (.A(_03529_),
    .B(_03534_),
    .Y(_03535_));
 sky130_fd_sc_hd__nand2_1 _09627_ (.A(_03535_),
    .B(_03274_),
    .Y(_03536_));
 sky130_fd_sc_hd__nand3_1 _09628_ (.A(_03230_),
    .B(_03406_),
    .C(_03231_),
    .Y(_03537_));
 sky130_fd_sc_hd__nand2_1 _09629_ (.A(_03403_),
    .B(_03381_),
    .Y(_03538_));
 sky130_fd_sc_hd__nor2_1 _09630_ (.A(_03381_),
    .B(_03403_),
    .Y(_03539_));
 sky130_fd_sc_hd__a21oi_1 _09631_ (.A1(_03538_),
    .A2(_03214_),
    .B1(_03539_),
    .Y(_03540_));
 sky130_fd_sc_hd__nand2_1 _09632_ (.A(_03537_),
    .B(_03540_),
    .Y(_03541_));
 sky130_fd_sc_hd__nor2_1 _09633_ (.A(_03507_),
    .B(_03206_),
    .Y(_03542_));
 sky130_fd_sc_hd__a21oi_1 _09634_ (.A1(_03389_),
    .A2(_03384_),
    .B1(_03386_),
    .Y(_03543_));
 sky130_fd_sc_hd__nor2_1 _09635_ (.A(_03350_),
    .B(_03383_),
    .Y(_03544_));
 sky130_fd_sc_hd__nand2_1 _09636_ (.A(_03076_),
    .B(_03020_),
    .Y(_03545_));
 sky130_fd_sc_hd__nand2_1 _09637_ (.A(_03110_),
    .B(_03020_),
    .Y(_03546_));
 sky130_fd_sc_hd__nand2_1 _09638_ (.A(_03385_),
    .B(_03546_),
    .Y(_03547_));
 sky130_fd_sc_hd__o21a_1 _09639_ (.A1(_03387_),
    .A2(_03545_),
    .B1(_03547_),
    .X(_03548_));
 sky130_fd_sc_hd__or2_1 _09640_ (.A(_03544_),
    .B(_03548_),
    .X(_03549_));
 sky130_fd_sc_hd__nand2_1 _09641_ (.A(_03548_),
    .B(_03544_),
    .Y(_03550_));
 sky130_fd_sc_hd__nand2_1 _09642_ (.A(_03549_),
    .B(_03550_),
    .Y(_03551_));
 sky130_fd_sc_hd__xor2_1 _09643_ (.A(_03543_),
    .B(_03551_),
    .X(_03552_));
 sky130_fd_sc_hd__nor2_1 _09644_ (.A(_03542_),
    .B(_03552_),
    .Y(_03553_));
 sky130_fd_sc_hd__nand2_1 _09645_ (.A(_03552_),
    .B(_03542_),
    .Y(_03554_));
 sky130_fd_sc_hd__inv_2 _09646_ (.A(_03554_),
    .Y(_03555_));
 sky130_fd_sc_hd__o21ai_1 _09647_ (.A1(_03395_),
    .A2(_03394_),
    .B1(_03401_),
    .Y(_03556_));
 sky130_fd_sc_hd__o21bai_1 _09648_ (.A1(_03553_),
    .A2(_03555_),
    .B1_N(_03556_),
    .Y(_03557_));
 sky130_fd_sc_hd__inv_2 _09649_ (.A(_03553_),
    .Y(_03558_));
 sky130_fd_sc_hd__nand3_1 _09650_ (.A(_03558_),
    .B(_03556_),
    .C(_03554_),
    .Y(_03559_));
 sky130_fd_sc_hd__nand2_1 _09651_ (.A(_03557_),
    .B(_03559_),
    .Y(_03560_));
 sky130_fd_sc_hd__inv_2 _09652_ (.A(_03560_),
    .Y(_03561_));
 sky130_fd_sc_hd__nand2_1 _09653_ (.A(_03541_),
    .B(_03561_),
    .Y(_03562_));
 sky130_fd_sc_hd__nand3_1 _09654_ (.A(_03560_),
    .B(_03537_),
    .C(_03540_),
    .Y(_03563_));
 sky130_fd_sc_hd__nand2_1 _09655_ (.A(_03562_),
    .B(_03563_),
    .Y(_03564_));
 sky130_fd_sc_hd__nand2_1 _09656_ (.A(_03564_),
    .B(_03233_),
    .Y(_03565_));
 sky130_fd_sc_hd__nand3_1 _09657_ (.A(_03536_),
    .B(_00623_),
    .C(_03565_),
    .Y(_03566_));
 sky130_fd_sc_hd__nand2_1 _09658_ (.A(_03110_),
    .B(_00556_),
    .Y(_03567_));
 sky130_fd_sc_hd__nand3_1 _09659_ (.A(_03566_),
    .B(_02092_),
    .C(_03567_),
    .Y(_03568_));
 sky130_fd_sc_hd__nand3_1 _09660_ (.A(_03529_),
    .B(_03534_),
    .C(_03274_),
    .Y(_03569_));
 sky130_fd_sc_hd__nand3_1 _09661_ (.A(_03562_),
    .B(_03563_),
    .C(_03233_),
    .Y(_03570_));
 sky130_fd_sc_hd__nand3_1 _09662_ (.A(_03569_),
    .B(_00623_),
    .C(_03570_),
    .Y(_03571_));
 sky130_fd_sc_hd__or2_1 _09663_ (.A(_00623_),
    .B(_03110_),
    .X(_03572_));
 sky130_fd_sc_hd__nand3_1 _09664_ (.A(_03571_),
    .B(_00831_),
    .C(_03572_),
    .Y(_03573_));
 sky130_fd_sc_hd__a21o_1 _09665_ (.A1(\H[3][6] ),
    .A2(_03033_),
    .B1(_03026_),
    .X(_03574_));
 sky130_fd_sc_hd__a21o_1 _09666_ (.A1(\H[2][6] ),
    .A2(_03022_),
    .B1(_03574_),
    .X(_03575_));
 sky130_fd_sc_hd__nor2_1 _09667_ (.A(_03025_),
    .B(_02303_),
    .Y(_03576_));
 sky130_fd_sc_hd__a211o_1 _09668_ (.A1(\H[1][6] ),
    .A2(_03025_),
    .B1(_02840_),
    .C1(_03576_),
    .X(_03577_));
 sky130_fd_sc_hd__nand2_1 _09669_ (.A(_03021_),
    .B(\Oset[0][6] ),
    .Y(_03578_));
 sky130_fd_sc_hd__nand2_1 _09670_ (.A(\Oset[1][6] ),
    .B(_03024_),
    .Y(_03579_));
 sky130_fd_sc_hd__a21oi_1 _09671_ (.A1(\Oset[3][6] ),
    .A2(_03024_),
    .B1(_03026_),
    .Y(_03580_));
 sky130_fd_sc_hd__nand2_1 _09672_ (.A(_03021_),
    .B(\Oset[2][6] ),
    .Y(_03581_));
 sky130_fd_sc_hd__a32o_1 _09673_ (.A1(_03578_),
    .A2(_03579_),
    .A3(_03026_),
    .B1(_03580_),
    .B2(_03581_),
    .X(_03582_));
 sky130_fd_sc_hd__nand2_1 _09674_ (.A(_03021_),
    .B(\Qset[0][6] ),
    .Y(_03583_));
 sky130_fd_sc_hd__nand2_1 _09675_ (.A(\Qset[1][6] ),
    .B(_03024_),
    .Y(_03584_));
 sky130_fd_sc_hd__a21oi_1 _09676_ (.A1(\Qset[3][6] ),
    .A2(_03024_),
    .B1(_03026_),
    .Y(_03585_));
 sky130_fd_sc_hd__nand2_1 _09677_ (.A(_03021_),
    .B(\Qset[2][6] ),
    .Y(_03586_));
 sky130_fd_sc_hd__a32o_1 _09678_ (.A1(_03583_),
    .A2(_03584_),
    .A3(_03026_),
    .B1(_03585_),
    .B2(_03586_),
    .X(_03587_));
 sky130_fd_sc_hd__mux2_1 _09679_ (.A0(_03582_),
    .A1(_03587_),
    .S(_00646_),
    .X(_03588_));
 sky130_fd_sc_hd__nor2_1 _09680_ (.A(_01536_),
    .B(_03588_),
    .Y(_03589_));
 sky130_fd_sc_hd__a311o_2 _09681_ (.A1(_01537_),
    .A2(_03575_),
    .A3(_03577_),
    .B1(_00549_),
    .C1(_03589_),
    .X(_03590_));
 sky130_fd_sc_hd__o21ai_2 _09682_ (.A1(_00623_),
    .A2(_03506_),
    .B1(_03590_),
    .Y(_03591_));
 sky130_fd_sc_hd__nand3_1 _09683_ (.A(_03568_),
    .B(_03573_),
    .C(_03591_),
    .Y(_03592_));
 sky130_fd_sc_hd__nand3_1 _09684_ (.A(_03566_),
    .B(_00536_),
    .C(_03567_),
    .Y(_03593_));
 sky130_fd_sc_hd__nand3_1 _09685_ (.A(_03571_),
    .B(_02092_),
    .C(_03572_),
    .Y(_03594_));
 sky130_fd_sc_hd__inv_2 _09686_ (.A(_03591_),
    .Y(_03595_));
 sky130_fd_sc_hd__nand3_1 _09687_ (.A(_03593_),
    .B(_03594_),
    .C(_03595_),
    .Y(_03596_));
 sky130_fd_sc_hd__nand2_1 _09688_ (.A(_03592_),
    .B(_03596_),
    .Y(_03597_));
 sky130_fd_sc_hd__nor2_1 _09689_ (.A(_03444_),
    .B(_03597_),
    .Y(_03598_));
 sky130_fd_sc_hd__and2_1 _09690_ (.A(_03597_),
    .B(_03444_),
    .X(_03599_));
 sky130_fd_sc_hd__or2_2 _09691_ (.A(_03598_),
    .B(_03599_),
    .X(_03600_));
 sky130_fd_sc_hd__xor2_4 _09692_ (.A(_03452_),
    .B(_03600_),
    .X(_03601_));
 sky130_fd_sc_hd__nor2_1 _09693_ (.A(_02653_),
    .B(_03601_),
    .Y(_03602_));
 sky130_fd_sc_hd__a211o_1 _09694_ (.A1(_00857_),
    .A2(_02654_),
    .B1(_02753_),
    .C1(_03602_),
    .X(_03603_));
 sky130_fd_sc_hd__inv_2 _09695_ (.A(_03603_),
    .Y(_00250_));
 sky130_fd_sc_hd__o21bai_2 _09696_ (.A1(_03452_),
    .A2(_03599_),
    .B1_N(_03598_),
    .Y(_03604_));
 sky130_fd_sc_hd__a21boi_1 _09697_ (.A1(_03528_),
    .A2(_03530_),
    .B1_N(_03531_),
    .Y(_03605_));
 sky130_fd_sc_hd__nor2_1 _09698_ (.A(_03514_),
    .B(_03511_),
    .Y(_03606_));
 sky130_fd_sc_hd__inv_2 _09699_ (.A(_03606_),
    .Y(_03607_));
 sky130_fd_sc_hd__nand2_1 _09700_ (.A(_03519_),
    .B(_03607_),
    .Y(_03608_));
 sky130_fd_sc_hd__nor2_1 _09701_ (.A(_03464_),
    .B(_03463_),
    .Y(_03609_));
 sky130_fd_sc_hd__a21oi_2 _09702_ (.A1(_03465_),
    .A2(_03461_),
    .B1(_03609_),
    .Y(_03610_));
 sky130_fd_sc_hd__inv_2 _09703_ (.A(_03610_),
    .Y(_03611_));
 sky130_fd_sc_hd__nand2_1 _09704_ (.A(_03421_),
    .B(_03462_),
    .Y(_03612_));
 sky130_fd_sc_hd__nand2_1 _09705_ (.A(_02895_),
    .B(_03079_),
    .Y(_03613_));
 sky130_fd_sc_hd__inv_2 _09706_ (.A(_03613_),
    .Y(_03614_));
 sky130_fd_sc_hd__nand3_1 _09707_ (.A(_03612_),
    .B(_03020_),
    .C(_03614_),
    .Y(_03615_));
 sky130_fd_sc_hd__nand2_1 _09708_ (.A(_03020_),
    .B(_03614_),
    .Y(_03616_));
 sky130_fd_sc_hd__nand3_1 _09709_ (.A(_03616_),
    .B(_03421_),
    .C(_03462_),
    .Y(_03617_));
 sky130_fd_sc_hd__nand2_1 _09710_ (.A(_03506_),
    .B(_03304_),
    .Y(_03618_));
 sky130_fd_sc_hd__nand3_1 _09711_ (.A(_03615_),
    .B(_03617_),
    .C(_03618_),
    .Y(_03619_));
 sky130_fd_sc_hd__a21oi_1 _09712_ (.A1(_03348_),
    .A2(_02286_),
    .B1(_03613_),
    .Y(_03620_));
 sky130_fd_sc_hd__nand2_1 _09713_ (.A(_03620_),
    .B(_03459_),
    .Y(_03621_));
 sky130_fd_sc_hd__a21oi_1 _09714_ (.A1(_03504_),
    .A2(_02308_),
    .B1(_03303_),
    .Y(_03622_));
 sky130_fd_sc_hd__nand2_1 _09715_ (.A(_03612_),
    .B(_03616_),
    .Y(_03623_));
 sky130_fd_sc_hd__nand3_2 _09716_ (.A(_03621_),
    .B(_03622_),
    .C(_03623_),
    .Y(_03624_));
 sky130_fd_sc_hd__nand3_1 _09717_ (.A(_03611_),
    .B(_03619_),
    .C(_03624_),
    .Y(_03625_));
 sky130_fd_sc_hd__nand2_1 _09718_ (.A(_03619_),
    .B(_03624_),
    .Y(_03626_));
 sky130_fd_sc_hd__nand2_1 _09719_ (.A(_03626_),
    .B(_03610_),
    .Y(_03627_));
 sky130_fd_sc_hd__nor2_1 _09720_ (.A(_03498_),
    .B(_02320_),
    .Y(_03628_));
 sky130_fd_sc_hd__a211o_1 _09721_ (.A1(_03498_),
    .A2(\Oset[3][7] ),
    .B1(_03004_),
    .C1(_03628_),
    .X(_03629_));
 sky130_fd_sc_hd__nor2_1 _09722_ (.A(_03498_),
    .B(_02323_),
    .Y(_03630_));
 sky130_fd_sc_hd__a211o_1 _09723_ (.A1(_03498_),
    .A2(\Oset[1][7] ),
    .B1(_02991_),
    .C1(_03630_),
    .X(_03631_));
 sky130_fd_sc_hd__nand2_2 _09724_ (.A(_03629_),
    .B(_03631_),
    .Y(_03632_));
 sky130_fd_sc_hd__o21ai_1 _09725_ (.A1(_02540_),
    .A2(_03632_),
    .B1(_01155_),
    .Y(_03633_));
 sky130_fd_sc_hd__nand2_1 _09726_ (.A(_02318_),
    .B(_02162_),
    .Y(_03634_));
 sky130_fd_sc_hd__nor2_1 _09727_ (.A(\Qset[3][7] ),
    .B(_03341_),
    .Y(_03635_));
 sky130_fd_sc_hd__o21ai_1 _09728_ (.A1(_02992_),
    .A2(\Qset[2][7] ),
    .B1(_02991_),
    .Y(_03636_));
 sky130_fd_sc_hd__nor2_1 _09729_ (.A(_03001_),
    .B(\Qset[0][7] ),
    .Y(_03637_));
 sky130_fd_sc_hd__o21ai_1 _09730_ (.A1(\Qset[1][7] ),
    .A2(_03341_),
    .B1(_03004_),
    .Y(_03638_));
 sky130_fd_sc_hd__o22a_2 _09731_ (.A1(_03635_),
    .A2(_03636_),
    .B1(_03637_),
    .B2(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__nand2_1 _09732_ (.A(_03639_),
    .B(_00581_),
    .Y(_03640_));
 sky130_fd_sc_hd__and3_1 _09733_ (.A(_03634_),
    .B(_03640_),
    .C(_02540_),
    .X(_03641_));
 sky130_fd_sc_hd__a21oi_1 _09734_ (.A1(_02326_),
    .A2(_00584_),
    .B1(_02573_),
    .Y(_03642_));
 sky130_fd_sc_hd__o21ai_1 _09735_ (.A1(_03633_),
    .A2(_03641_),
    .B1(_03642_),
    .Y(_03643_));
 sky130_fd_sc_hd__mux2_1 _09736_ (.A0(\H[2][7] ),
    .A1(\H[3][7] ),
    .S(_02611_),
    .X(_03644_));
 sky130_fd_sc_hd__nor2_1 _09737_ (.A(_03498_),
    .B(\H[0][7] ),
    .Y(_03645_));
 sky130_fd_sc_hd__o21ai_1 _09738_ (.A1(\H[1][7] ),
    .A2(_03341_),
    .B1(_03004_),
    .Y(_03646_));
 sky130_fd_sc_hd__o2bb2a_1 _09739_ (.A1_N(_02991_),
    .A2_N(_03644_),
    .B1(_03645_),
    .B2(_03646_),
    .X(_03647_));
 sky130_fd_sc_hd__or2_1 _09740_ (.A(_02556_),
    .B(_03647_),
    .X(_03648_));
 sky130_fd_sc_hd__nand2_1 _09741_ (.A(_03643_),
    .B(_03648_),
    .Y(_03649_));
 sky130_fd_sc_hd__nand2_1 _09742_ (.A(_03649_),
    .B(_01552_),
    .Y(_03650_));
 sky130_fd_sc_hd__nand2_4 _09743_ (.A(_03650_),
    .B(_02334_),
    .Y(_03651_));
 sky130_fd_sc_hd__buf_6 _09744_ (.A(_03651_),
    .X(_03652_));
 sky130_fd_sc_hd__nand2_1 _09745_ (.A(_03652_),
    .B(_03257_),
    .Y(_03653_));
 sky130_fd_sc_hd__inv_2 _09746_ (.A(_03653_),
    .Y(_03654_));
 sky130_fd_sc_hd__nand3_1 _09747_ (.A(_03625_),
    .B(_03627_),
    .C(_03654_),
    .Y(_03655_));
 sky130_fd_sc_hd__nand2_1 _09748_ (.A(_03626_),
    .B(_03611_),
    .Y(_03656_));
 sky130_fd_sc_hd__nand3_1 _09749_ (.A(_03619_),
    .B(_03624_),
    .C(_03610_),
    .Y(_03657_));
 sky130_fd_sc_hd__nand3_1 _09750_ (.A(_03656_),
    .B(_03657_),
    .C(_03653_),
    .Y(_03658_));
 sky130_fd_sc_hd__nand2_1 _09751_ (.A(_03655_),
    .B(_03658_),
    .Y(_03659_));
 sky130_fd_sc_hd__nand2_1 _09752_ (.A(_03471_),
    .B(_03473_),
    .Y(_03660_));
 sky130_fd_sc_hd__nor2_1 _09753_ (.A(_03473_),
    .B(_03471_),
    .Y(_03661_));
 sky130_fd_sc_hd__a21oi_1 _09754_ (.A1(_03660_),
    .A2(_03508_),
    .B1(_03661_),
    .Y(_03662_));
 sky130_fd_sc_hd__inv_2 _09755_ (.A(_03662_),
    .Y(_03663_));
 sky130_fd_sc_hd__nand2_1 _09756_ (.A(_03659_),
    .B(_03663_),
    .Y(_03664_));
 sky130_fd_sc_hd__nand3_1 _09757_ (.A(_03662_),
    .B(_03655_),
    .C(_03658_),
    .Y(_03665_));
 sky130_fd_sc_hd__nand2_1 _09758_ (.A(_03664_),
    .B(_03665_),
    .Y(_03666_));
 sky130_fd_sc_hd__nand2_1 _09759_ (.A(_03608_),
    .B(_03666_),
    .Y(_03667_));
 sky130_fd_sc_hd__nand3b_1 _09760_ (.A_N(_03666_),
    .B(_03519_),
    .C(_03607_),
    .Y(_03668_));
 sky130_fd_sc_hd__nand2_1 _09761_ (.A(_03667_),
    .B(_03668_),
    .Y(_03669_));
 sky130_fd_sc_hd__a21o_1 _09762_ (.A1(_03218_),
    .A2(_03219_),
    .B1(_03227_),
    .X(_03670_));
 sky130_fd_sc_hd__nand2_1 _09763_ (.A(_03670_),
    .B(_03228_),
    .Y(_03671_));
 sky130_fd_sc_hd__nand2_1 _09764_ (.A(_03669_),
    .B(_03671_),
    .Y(_03672_));
 sky130_fd_sc_hd__inv_2 _09765_ (.A(_03671_),
    .Y(_03673_));
 sky130_fd_sc_hd__nand3_1 _09766_ (.A(_03667_),
    .B(_03668_),
    .C(_03673_),
    .Y(_03674_));
 sky130_fd_sc_hd__nand2_1 _09767_ (.A(_03672_),
    .B(_03674_),
    .Y(_03675_));
 sky130_fd_sc_hd__nand2_1 _09768_ (.A(_03605_),
    .B(_03675_),
    .Y(_03676_));
 sky130_fd_sc_hd__nand2_1 _09769_ (.A(_03529_),
    .B(_03531_),
    .Y(_03677_));
 sky130_fd_sc_hd__nand2_1 _09770_ (.A(_03669_),
    .B(_03673_),
    .Y(_03678_));
 sky130_fd_sc_hd__nand3_1 _09771_ (.A(_03667_),
    .B(_03668_),
    .C(_03671_),
    .Y(_03679_));
 sky130_fd_sc_hd__nand2_1 _09772_ (.A(_03678_),
    .B(_03679_),
    .Y(_03680_));
 sky130_fd_sc_hd__nand2_1 _09773_ (.A(_03677_),
    .B(_03680_),
    .Y(_03681_));
 sky130_fd_sc_hd__nand3_1 _09774_ (.A(_03676_),
    .B(_03681_),
    .C(_03274_),
    .Y(_03682_));
 sky130_fd_sc_hd__nand2_1 _09775_ (.A(_03562_),
    .B(_03559_),
    .Y(_03683_));
 sky130_fd_sc_hd__o21a_1 _09776_ (.A1(_03543_),
    .A2(_03551_),
    .B1(_03554_),
    .X(_03684_));
 sky130_fd_sc_hd__inv_2 _09777_ (.A(_03651_),
    .Y(_03685_));
 sky130_fd_sc_hd__nor2_1 _09778_ (.A(_03206_),
    .B(_03685_),
    .Y(_03686_));
 sky130_fd_sc_hd__nor2_1 _09779_ (.A(_03507_),
    .B(_03383_),
    .Y(_03687_));
 sky130_fd_sc_hd__nand2_1 _09780_ (.A(_03076_),
    .B(_03421_),
    .Y(_03688_));
 sky130_fd_sc_hd__or2_1 _09781_ (.A(_03546_),
    .B(_03688_),
    .X(_03689_));
 sky130_fd_sc_hd__nand2_1 _09782_ (.A(_03110_),
    .B(_03421_),
    .Y(_03690_));
 sky130_fd_sc_hd__nand2_1 _09783_ (.A(_03545_),
    .B(_03690_),
    .Y(_03691_));
 sky130_fd_sc_hd__nand2_1 _09784_ (.A(_03689_),
    .B(_03691_),
    .Y(_03692_));
 sky130_fd_sc_hd__xor2_1 _09785_ (.A(_03687_),
    .B(_03692_),
    .X(_03693_));
 sky130_fd_sc_hd__o21a_1 _09786_ (.A1(_03385_),
    .A2(_03546_),
    .B1(_03550_),
    .X(_03694_));
 sky130_fd_sc_hd__or2_1 _09787_ (.A(_03693_),
    .B(_03694_),
    .X(_03695_));
 sky130_fd_sc_hd__nand2_1 _09788_ (.A(_03694_),
    .B(_03693_),
    .Y(_03696_));
 sky130_fd_sc_hd__nand2_1 _09789_ (.A(_03695_),
    .B(_03696_),
    .Y(_03697_));
 sky130_fd_sc_hd__xor2_1 _09790_ (.A(_03686_),
    .B(_03697_),
    .X(_03698_));
 sky130_fd_sc_hd__or2_1 _09791_ (.A(_03684_),
    .B(_03698_),
    .X(_03699_));
 sky130_fd_sc_hd__nand2_1 _09792_ (.A(_03698_),
    .B(_03684_),
    .Y(_03700_));
 sky130_fd_sc_hd__nand3_1 _09793_ (.A(_03683_),
    .B(_03699_),
    .C(_03700_),
    .Y(_03701_));
 sky130_fd_sc_hd__nand2_1 _09794_ (.A(_03699_),
    .B(_03700_),
    .Y(_03702_));
 sky130_fd_sc_hd__nand3_1 _09795_ (.A(_03562_),
    .B(_03702_),
    .C(_03559_),
    .Y(_03703_));
 sky130_fd_sc_hd__nand3_2 _09796_ (.A(_03701_),
    .B(_03703_),
    .C(_03233_),
    .Y(_03704_));
 sky130_fd_sc_hd__nand3_1 _09797_ (.A(_03682_),
    .B(_03704_),
    .C(_00624_),
    .Y(_03705_));
 sky130_fd_sc_hd__or2_1 _09798_ (.A(_00623_),
    .B(_03076_),
    .X(_03706_));
 sky130_fd_sc_hd__nand2_1 _09799_ (.A(_03705_),
    .B(_03706_),
    .Y(_03707_));
 sky130_fd_sc_hd__nand2_1 _09800_ (.A(_03707_),
    .B(_00831_),
    .Y(_03708_));
 sky130_fd_sc_hd__nand3_1 _09801_ (.A(_03705_),
    .B(_02092_),
    .C(_03706_),
    .Y(_03709_));
 sky130_fd_sc_hd__a21o_1 _09802_ (.A1(\H[3][7] ),
    .A2(_03025_),
    .B1(_03027_),
    .X(_03710_));
 sky130_fd_sc_hd__a21o_1 _09803_ (.A1(\H[2][7] ),
    .A2(_03023_),
    .B1(_03710_),
    .X(_03711_));
 sky130_fd_sc_hd__a21o_1 _09804_ (.A1(\H[1][7] ),
    .A2(_03025_),
    .B1(_02840_),
    .X(_03712_));
 sky130_fd_sc_hd__a21o_1 _09805_ (.A1(\H[0][7] ),
    .A2(_03022_),
    .B1(_03712_),
    .X(_03713_));
 sky130_fd_sc_hd__nand2_1 _09806_ (.A(_03021_),
    .B(\Oset[0][7] ),
    .Y(_03714_));
 sky130_fd_sc_hd__nand2_1 _09807_ (.A(\Oset[1][7] ),
    .B(_03033_),
    .Y(_03715_));
 sky130_fd_sc_hd__a21oi_1 _09808_ (.A1(\Oset[3][7] ),
    .A2(_03033_),
    .B1(_03026_),
    .Y(_03716_));
 sky130_fd_sc_hd__nand2_1 _09809_ (.A(_03022_),
    .B(\Oset[2][7] ),
    .Y(_03717_));
 sky130_fd_sc_hd__a32o_1 _09810_ (.A1(_03714_),
    .A2(_03715_),
    .A3(_03027_),
    .B1(_03716_),
    .B2(_03717_),
    .X(_03718_));
 sky130_fd_sc_hd__nand2_1 _09811_ (.A(_03021_),
    .B(\Qset[0][7] ),
    .Y(_03719_));
 sky130_fd_sc_hd__nand2_1 _09812_ (.A(\Qset[1][7] ),
    .B(_03033_),
    .Y(_03720_));
 sky130_fd_sc_hd__a21oi_1 _09813_ (.A1(\Qset[3][7] ),
    .A2(_03033_),
    .B1(_03026_),
    .Y(_03721_));
 sky130_fd_sc_hd__nand2_1 _09814_ (.A(_03022_),
    .B(\Qset[2][7] ),
    .Y(_03722_));
 sky130_fd_sc_hd__a32o_1 _09815_ (.A1(_03719_),
    .A2(_03720_),
    .A3(_03027_),
    .B1(_03721_),
    .B2(_03722_),
    .X(_03723_));
 sky130_fd_sc_hd__mux2_1 _09816_ (.A0(_03718_),
    .A1(_03723_),
    .S(_00647_),
    .X(_03724_));
 sky130_fd_sc_hd__nor2_1 _09817_ (.A(_01537_),
    .B(_03724_),
    .Y(_03725_));
 sky130_fd_sc_hd__a311o_2 _09818_ (.A1(_01537_),
    .A2(_03711_),
    .A3(_03713_),
    .B1(_00549_),
    .C1(_03725_),
    .X(_03726_));
 sky130_fd_sc_hd__o21ai_2 _09819_ (.A1(_00624_),
    .A2(_03652_),
    .B1(_03726_),
    .Y(_03727_));
 sky130_fd_sc_hd__inv_2 _09820_ (.A(_03727_),
    .Y(_03728_));
 sky130_fd_sc_hd__nand3_1 _09821_ (.A(_03708_),
    .B(_03709_),
    .C(_03728_),
    .Y(_03729_));
 sky130_fd_sc_hd__nand2_1 _09822_ (.A(_03707_),
    .B(_02092_),
    .Y(_03730_));
 sky130_fd_sc_hd__nand3_1 _09823_ (.A(_03705_),
    .B(_00831_),
    .C(_03706_),
    .Y(_03731_));
 sky130_fd_sc_hd__nand3_1 _09824_ (.A(_03730_),
    .B(_03731_),
    .C(_03727_),
    .Y(_03732_));
 sky130_fd_sc_hd__nand2_1 _09825_ (.A(_03729_),
    .B(_03732_),
    .Y(_03733_));
 sky130_fd_sc_hd__inv_2 _09826_ (.A(_03596_),
    .Y(_03734_));
 sky130_fd_sc_hd__nand2_1 _09827_ (.A(_03733_),
    .B(_03734_),
    .Y(_03735_));
 sky130_fd_sc_hd__nand3_1 _09828_ (.A(_03729_),
    .B(_03732_),
    .C(_03596_),
    .Y(_03736_));
 sky130_fd_sc_hd__nand2_1 _09829_ (.A(_03735_),
    .B(_03736_),
    .Y(_03737_));
 sky130_fd_sc_hd__or2_1 _09830_ (.A(_03604_),
    .B(_03737_),
    .X(_03738_));
 sky130_fd_sc_hd__nand2_1 _09831_ (.A(_03737_),
    .B(_03604_),
    .Y(_03739_));
 sky130_fd_sc_hd__and2_2 _09832_ (.A(_03738_),
    .B(_03739_),
    .X(_03740_));
 sky130_fd_sc_hd__nor2_1 _09833_ (.A(_02653_),
    .B(_03740_),
    .Y(_03741_));
 sky130_fd_sc_hd__a211o_1 _09834_ (.A1(_00884_),
    .A2(_02654_),
    .B1(_02753_),
    .C1(_03741_),
    .X(_03742_));
 sky130_fd_sc_hd__inv_2 _09835_ (.A(_03742_),
    .Y(_00251_));
 sky130_fd_sc_hd__inv_2 _09836_ (.A(_03729_),
    .Y(_03743_));
 sky130_fd_sc_hd__nand3_1 _09837_ (.A(_03604_),
    .B(_03734_),
    .C(_03743_),
    .Y(_03744_));
 sky130_fd_sc_hd__clkbuf_4 _09838_ (.A(_03050_),
    .X(_03745_));
 sky130_fd_sc_hd__buf_6 _09839_ (.A(_03745_),
    .X(_03746_));
 sky130_fd_sc_hd__nand2_1 _09840_ (.A(_03744_),
    .B(_03746_),
    .Y(_03747_));
 sky130_fd_sc_hd__inv_2 _09841_ (.A(_03747_),
    .Y(_03748_));
 sky130_fd_sc_hd__a21oi_1 _09842_ (.A1(_03732_),
    .A2(_03734_),
    .B1(_03743_),
    .Y(_03749_));
 sky130_fd_sc_hd__nand2_1 _09843_ (.A(_03739_),
    .B(_03749_),
    .Y(_03750_));
 sky130_fd_sc_hd__buf_4 _09844_ (.A(_03047_),
    .X(_03751_));
 sky130_fd_sc_hd__a21o_1 _09845_ (.A1(_03280_),
    .A2(_03751_),
    .B1(_00831_),
    .X(_03752_));
 sky130_fd_sc_hd__inv_2 _09846_ (.A(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__nand3_1 _09847_ (.A(_03748_),
    .B(_03750_),
    .C(_03753_),
    .Y(_03754_));
 sky130_fd_sc_hd__nand3_1 _09848_ (.A(_03750_),
    .B(_03746_),
    .C(_03744_),
    .Y(_03755_));
 sky130_fd_sc_hd__nand2_1 _09849_ (.A(_03755_),
    .B(_03752_),
    .Y(_03756_));
 sky130_fd_sc_hd__nand2_1 _09850_ (.A(_03754_),
    .B(_03756_),
    .Y(_03757_));
 sky130_fd_sc_hd__buf_4 _09851_ (.A(_02556_),
    .X(_03758_));
 sky130_fd_sc_hd__buf_6 _09852_ (.A(_03498_),
    .X(_03759_));
 sky130_fd_sc_hd__buf_6 _09853_ (.A(_03759_),
    .X(_03760_));
 sky130_fd_sc_hd__clkbuf_4 _09854_ (.A(_03004_),
    .X(_03761_));
 sky130_fd_sc_hd__nor2_1 _09855_ (.A(_03760_),
    .B(_02346_),
    .Y(_03762_));
 sky130_fd_sc_hd__a211o_1 _09856_ (.A1(_03760_),
    .A2(\H[3][8] ),
    .B1(_03761_),
    .C1(_03762_),
    .X(_03763_));
 sky130_fd_sc_hd__clkbuf_4 _09857_ (.A(_03345_),
    .X(_03764_));
 sky130_fd_sc_hd__nor2_1 _09858_ (.A(_03760_),
    .B(_02350_),
    .Y(_03765_));
 sky130_fd_sc_hd__a211o_1 _09859_ (.A1(_03760_),
    .A2(\H[1][8] ),
    .B1(_03764_),
    .C1(_03765_),
    .X(_03766_));
 sky130_fd_sc_hd__nand2_2 _09860_ (.A(_03763_),
    .B(_03766_),
    .Y(_03767_));
 sky130_fd_sc_hd__buf_4 _09861_ (.A(_02573_),
    .X(_03768_));
 sky130_fd_sc_hd__a21o_1 _09862_ (.A1(_02345_),
    .A2(_00584_),
    .B1(_03768_),
    .X(_03769_));
 sky130_fd_sc_hd__buf_4 _09863_ (.A(_02540_),
    .X(_03770_));
 sky130_fd_sc_hd__mux2_1 _09864_ (.A0(\Oset[2][8] ),
    .A1(\Oset[3][8] ),
    .S(_03498_),
    .X(_03771_));
 sky130_fd_sc_hd__nor2_1 _09865_ (.A(_03759_),
    .B(\Oset[0][8] ),
    .Y(_03772_));
 sky130_fd_sc_hd__buf_6 _09866_ (.A(_03341_),
    .X(_03773_));
 sky130_fd_sc_hd__o21ai_1 _09867_ (.A1(\Oset[1][8] ),
    .A2(_03773_),
    .B1(_03761_),
    .Y(_03774_));
 sky130_fd_sc_hd__o2bb2a_2 _09868_ (.A1_N(_03345_),
    .A2_N(_03771_),
    .B1(_03772_),
    .B2(_03774_),
    .X(_03775_));
 sky130_fd_sc_hd__nor2_1 _09869_ (.A(\Qset[3][8] ),
    .B(_03341_),
    .Y(_03776_));
 sky130_fd_sc_hd__o21ai_1 _09870_ (.A1(_03759_),
    .A2(\Qset[2][8] ),
    .B1(_03345_),
    .Y(_03777_));
 sky130_fd_sc_hd__nor2_1 _09871_ (.A(_03759_),
    .B(\Qset[0][8] ),
    .Y(_03778_));
 sky130_fd_sc_hd__o21ai_1 _09872_ (.A1(\Qset[1][8] ),
    .A2(_03773_),
    .B1(_03004_),
    .Y(_03779_));
 sky130_fd_sc_hd__o22a_2 _09873_ (.A1(_03776_),
    .A2(_03777_),
    .B1(_03778_),
    .B2(_03779_),
    .X(_03780_));
 sky130_fd_sc_hd__clkbuf_4 _09874_ (.A(_02552_),
    .X(_03781_));
 sky130_fd_sc_hd__a21oi_1 _09875_ (.A1(_03780_),
    .A2(_00582_),
    .B1(_03781_),
    .Y(_03782_));
 sky130_fd_sc_hd__nand2_1 _09876_ (.A(_02341_),
    .B(_02162_),
    .Y(_03783_));
 sky130_fd_sc_hd__nand2_1 _09877_ (.A(_03782_),
    .B(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__o21ai_1 _09878_ (.A1(_03770_),
    .A2(_03775_),
    .B1(_03784_),
    .Y(_03785_));
 sky130_fd_sc_hd__nor2_1 _09879_ (.A(_00584_),
    .B(_03785_),
    .Y(_03786_));
 sky130_fd_sc_hd__o22ai_1 _09880_ (.A1(_03758_),
    .A2(_03767_),
    .B1(_03769_),
    .B2(_03786_),
    .Y(_03787_));
 sky130_fd_sc_hd__nand2_1 _09881_ (.A(_03787_),
    .B(_01553_),
    .Y(_03788_));
 sky130_fd_sc_hd__nand2_2 _09882_ (.A(_03788_),
    .B(_02353_),
    .Y(_03789_));
 sky130_fd_sc_hd__buf_6 _09883_ (.A(_03789_),
    .X(_03790_));
 sky130_fd_sc_hd__clkbuf_4 _09884_ (.A(_03025_),
    .X(_03791_));
 sky130_fd_sc_hd__clkbuf_4 _09885_ (.A(_03791_),
    .X(_03792_));
 sky130_fd_sc_hd__buf_4 _09886_ (.A(_03792_),
    .X(_03793_));
 sky130_fd_sc_hd__clkbuf_4 _09887_ (.A(_03027_),
    .X(_03794_));
 sky130_fd_sc_hd__clkbuf_4 _09888_ (.A(_03794_),
    .X(_03795_));
 sky130_fd_sc_hd__nor2_1 _09889_ (.A(_03793_),
    .B(_02346_),
    .Y(_03796_));
 sky130_fd_sc_hd__a211o_1 _09890_ (.A1(\H[3][8] ),
    .A2(_03793_),
    .B1(_03795_),
    .C1(_03796_),
    .X(_03797_));
 sky130_fd_sc_hd__clkbuf_4 _09891_ (.A(_02840_),
    .X(_03798_));
 sky130_fd_sc_hd__nor2_1 _09892_ (.A(_03792_),
    .B(_02350_),
    .Y(_03799_));
 sky130_fd_sc_hd__a211o_1 _09893_ (.A1(\H[1][8] ),
    .A2(_03793_),
    .B1(_03798_),
    .C1(_03799_),
    .X(_03800_));
 sky130_fd_sc_hd__mux2_1 _09894_ (.A0(\Oset[0][8] ),
    .A1(\Oset[1][8] ),
    .S(_03791_),
    .X(_03801_));
 sky130_fd_sc_hd__or2_1 _09895_ (.A(\Oset[2][8] ),
    .B(_03791_),
    .X(_03802_));
 sky130_fd_sc_hd__o211a_1 _09896_ (.A1(\Oset[3][8] ),
    .A2(_03023_),
    .B1(_03798_),
    .C1(_03802_),
    .X(_03803_));
 sky130_fd_sc_hd__a211o_1 _09897_ (.A1(_03801_),
    .A2(_03794_),
    .B1(_00647_),
    .C1(_03803_),
    .X(_03804_));
 sky130_fd_sc_hd__mux2_1 _09898_ (.A0(\Qset[0][8] ),
    .A1(\Qset[1][8] ),
    .S(_03791_),
    .X(_03805_));
 sky130_fd_sc_hd__or2_1 _09899_ (.A(\Qset[2][8] ),
    .B(_03025_),
    .X(_03806_));
 sky130_fd_sc_hd__o211a_1 _09900_ (.A1(\Qset[3][8] ),
    .A2(_03023_),
    .B1(_03798_),
    .C1(_03806_),
    .X(_03807_));
 sky130_fd_sc_hd__a211o_1 _09901_ (.A1(_03805_),
    .A2(_03794_),
    .B1(_00621_),
    .C1(_03807_),
    .X(_03808_));
 sky130_fd_sc_hd__a31o_1 _09902_ (.A1(_03804_),
    .A2(_03808_),
    .A3(_00626_),
    .B1(_00556_),
    .X(_03809_));
 sky130_fd_sc_hd__a31o_2 _09903_ (.A1(_01538_),
    .A2(_03797_),
    .A3(_03800_),
    .B1(_03809_),
    .X(_03810_));
 sky130_fd_sc_hd__o21ai_2 _09904_ (.A1(_00624_),
    .A2(_03790_),
    .B1(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hd__nand2_1 _09905_ (.A(_03757_),
    .B(_03811_),
    .Y(_03812_));
 sky130_fd_sc_hd__inv_2 _09906_ (.A(_03811_),
    .Y(_03813_));
 sky130_fd_sc_hd__nand3_1 _09907_ (.A(_03754_),
    .B(_03756_),
    .C(_03813_),
    .Y(_03814_));
 sky130_fd_sc_hd__nor2_1 _09908_ (.A(\Qset[3][8] ),
    .B(_03136_),
    .Y(_03815_));
 sky130_fd_sc_hd__o21ai_1 _09909_ (.A1(_02545_),
    .A2(\Qset[2][8] ),
    .B1(_02526_),
    .Y(_03816_));
 sky130_fd_sc_hd__nor2_1 _09910_ (.A(_03157_),
    .B(\Qset[0][8] ),
    .Y(_03817_));
 sky130_fd_sc_hd__o21ai_1 _09911_ (.A1(\Qset[1][8] ),
    .A2(_03136_),
    .B1(_03135_),
    .Y(_03818_));
 sky130_fd_sc_hd__o22a_2 _09912_ (.A1(_03815_),
    .A2(_03816_),
    .B1(_03817_),
    .B2(_03818_),
    .X(_03819_));
 sky130_fd_sc_hd__o21ai_1 _09913_ (.A1(_02162_),
    .A2(_03819_),
    .B1(_02542_),
    .Y(_03820_));
 sky130_fd_sc_hd__or2_1 _09914_ (.A(_02562_),
    .B(\Oset[0][8] ),
    .X(_03821_));
 sky130_fd_sc_hd__o21a_1 _09915_ (.A1(\Oset[1][8] ),
    .A2(_02523_),
    .B1(_02535_),
    .X(_03822_));
 sky130_fd_sc_hd__mux2_1 _09916_ (.A0(\Oset[2][8] ),
    .A1(\Oset[3][8] ),
    .S(_02798_),
    .X(_03823_));
 sky130_fd_sc_hd__a22oi_4 _09917_ (.A1(_03821_),
    .A2(_03822_),
    .B1(_03823_),
    .B2(_02560_),
    .Y(_03824_));
 sky130_fd_sc_hd__nand2_1 _09918_ (.A(_03824_),
    .B(_02552_),
    .Y(_03825_));
 sky130_fd_sc_hd__nand3_1 _09919_ (.A(_03820_),
    .B(_03825_),
    .C(_01155_),
    .Y(_03826_));
 sky130_fd_sc_hd__nand2_1 _09920_ (.A(_03826_),
    .B(_02558_),
    .Y(_03827_));
 sky130_fd_sc_hd__mux2_1 _09921_ (.A0(\H[2][8] ),
    .A1(\H[3][8] ),
    .S(_02529_),
    .X(_03828_));
 sky130_fd_sc_hd__nor2_1 _09922_ (.A(_02565_),
    .B(_02350_),
    .Y(_03829_));
 sky130_fd_sc_hd__a211o_1 _09923_ (.A1(_02567_),
    .A2(\H[1][8] ),
    .B1(_02560_),
    .C1(_03829_),
    .X(_03830_));
 sky130_fd_sc_hd__o21ai_4 _09924_ (.A1(_03135_),
    .A2(_03828_),
    .B1(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__a21oi_1 _09925_ (.A1(_03831_),
    .A2(_02573_),
    .B1(_00588_),
    .Y(_03832_));
 sky130_fd_sc_hd__nand2_1 _09926_ (.A(_03827_),
    .B(_03832_),
    .Y(_03833_));
 sky130_fd_sc_hd__nand2_1 _09927_ (.A(_00588_),
    .B(\im_reg[8] ),
    .Y(_03834_));
 sky130_fd_sc_hd__nand2_4 _09928_ (.A(_03833_),
    .B(_03834_),
    .Y(_03835_));
 sky130_fd_sc_hd__nor2_1 _09929_ (.A(\Qset[3][9] ),
    .B(_03136_),
    .Y(_03836_));
 sky130_fd_sc_hd__o21ai_1 _09930_ (.A1(_03157_),
    .A2(\Qset[2][9] ),
    .B1(_02526_),
    .Y(_03837_));
 sky130_fd_sc_hd__nor2_1 _09931_ (.A(_02565_),
    .B(\Qset[0][9] ),
    .Y(_03838_));
 sky130_fd_sc_hd__o21ai_1 _09932_ (.A1(\Qset[1][9] ),
    .A2(_03136_),
    .B1(_03135_),
    .Y(_03839_));
 sky130_fd_sc_hd__o22a_4 _09933_ (.A1(_03836_),
    .A2(_03837_),
    .B1(_03838_),
    .B2(_03839_),
    .X(_03840_));
 sky130_fd_sc_hd__o21ai_1 _09934_ (.A1(_02162_),
    .A2(_03840_),
    .B1(_02713_),
    .Y(_03841_));
 sky130_fd_sc_hd__nor2_1 _09935_ (.A(_03157_),
    .B(_02368_),
    .Y(_03842_));
 sky130_fd_sc_hd__a211o_1 _09936_ (.A1(_02565_),
    .A2(\Oset[1][9] ),
    .B1(_02526_),
    .C1(_03842_),
    .X(_03843_));
 sky130_fd_sc_hd__nor2_1 _09937_ (.A(_02545_),
    .B(_02365_),
    .Y(_03844_));
 sky130_fd_sc_hd__a211o_1 _09938_ (.A1(_03157_),
    .A2(\Oset[3][9] ),
    .B1(_03135_),
    .C1(_03844_),
    .X(_03845_));
 sky130_fd_sc_hd__nand2_2 _09939_ (.A(_03843_),
    .B(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__nand2_1 _09940_ (.A(_03846_),
    .B(_03781_),
    .Y(_03847_));
 sky130_fd_sc_hd__nand3_1 _09941_ (.A(_03841_),
    .B(_01156_),
    .C(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__nand2_1 _09942_ (.A(_03848_),
    .B(_02723_),
    .Y(_03849_));
 sky130_fd_sc_hd__nor2_1 _09943_ (.A(_02567_),
    .B(\H[0][9] ),
    .Y(_03850_));
 sky130_fd_sc_hd__nor2_1 _09944_ (.A(\H[1][9] ),
    .B(_03152_),
    .Y(_03851_));
 sky130_fd_sc_hd__nor2_1 _09945_ (.A(_02565_),
    .B(\H[2][9] ),
    .Y(_03852_));
 sky130_fd_sc_hd__a211o_1 _09946_ (.A1(_02372_),
    .A2(_02565_),
    .B1(_03135_),
    .C1(_03852_),
    .X(_03853_));
 sky130_fd_sc_hd__o31a_2 _09947_ (.A1(_02560_),
    .A2(_03850_),
    .A3(_03851_),
    .B1(_03853_),
    .X(_03854_));
 sky130_fd_sc_hd__a21oi_1 _09948_ (.A1(_03854_),
    .A2(_02573_),
    .B1(_00588_),
    .Y(_03855_));
 sky130_fd_sc_hd__nand2_1 _09949_ (.A(_03849_),
    .B(_03855_),
    .Y(_03856_));
 sky130_fd_sc_hd__nand2_1 _09950_ (.A(_00588_),
    .B(\im_reg[9] ),
    .Y(_03857_));
 sky130_fd_sc_hd__nand2_2 _09951_ (.A(_03856_),
    .B(_03857_),
    .Y(_03858_));
 sky130_fd_sc_hd__buf_6 _09952_ (.A(_03858_),
    .X(_03859_));
 sky130_fd_sc_hd__nand3_1 _09953_ (.A(_03859_),
    .B(_02963_),
    .C(_03745_),
    .Y(_03860_));
 sky130_fd_sc_hd__inv_2 _09954_ (.A(\H[0][11] ),
    .Y(_03861_));
 sky130_fd_sc_hd__nand2_1 _09955_ (.A(_02787_),
    .B(_03861_),
    .Y(_03862_));
 sky130_fd_sc_hd__nand2_1 _09956_ (.A(_02423_),
    .B(_02528_),
    .Y(_03863_));
 sky130_fd_sc_hd__o21a_1 _09957_ (.A1(_02561_),
    .A2(\H[2][11] ),
    .B1(_02727_),
    .X(_03864_));
 sky130_fd_sc_hd__nand2_1 _09958_ (.A(_02420_),
    .B(_02544_),
    .Y(_03865_));
 sky130_fd_sc_hd__a32o_2 _09959_ (.A1(_03862_),
    .A2(_03863_),
    .A3(_02800_),
    .B1(_03864_),
    .B2(_03865_),
    .X(_03866_));
 sky130_fd_sc_hd__and3_1 _09960_ (.A(_03866_),
    .B(_01552_),
    .C(_02572_),
    .X(_03867_));
 sky130_fd_sc_hd__buf_4 _09961_ (.A(_03867_),
    .X(_03868_));
 sky130_fd_sc_hd__nand2_1 _09962_ (.A(_02785_),
    .B(_03868_),
    .Y(_03869_));
 sky130_fd_sc_hd__or2_1 _09963_ (.A(_02527_),
    .B(\H[0][10] ),
    .X(_03870_));
 sky130_fd_sc_hd__nand2_1 _09964_ (.A(_02400_),
    .B(_02874_),
    .Y(_03871_));
 sky130_fd_sc_hd__o21a_1 _09965_ (.A1(_02561_),
    .A2(\H[2][10] ),
    .B1(_02727_),
    .X(_03872_));
 sky130_fd_sc_hd__nand2_1 _09966_ (.A(_02396_),
    .B(_02544_),
    .Y(_03873_));
 sky130_fd_sc_hd__a32o_2 _09967_ (.A1(_03870_),
    .A2(_03871_),
    .A3(_02800_),
    .B1(_03872_),
    .B2(_03873_),
    .X(_03874_));
 sky130_fd_sc_hd__and3_1 _09968_ (.A(_03874_),
    .B(_01552_),
    .C(_02572_),
    .X(_03875_));
 sky130_fd_sc_hd__buf_4 _09969_ (.A(_03875_),
    .X(_03876_));
 sky130_fd_sc_hd__nand2_1 _09970_ (.A(_02687_),
    .B(_03876_),
    .Y(_03877_));
 sky130_fd_sc_hd__or2_1 _09971_ (.A(_03869_),
    .B(_03877_),
    .X(_03878_));
 sky130_fd_sc_hd__nand2_1 _09972_ (.A(_02784_),
    .B(_03876_),
    .Y(_03879_));
 sky130_fd_sc_hd__nand2_1 _09973_ (.A(_02687_),
    .B(_03868_),
    .Y(_03880_));
 sky130_fd_sc_hd__nand2_1 _09974_ (.A(_03879_),
    .B(_03880_),
    .Y(_03881_));
 sky130_fd_sc_hd__nand2_1 _09975_ (.A(_03878_),
    .B(_03881_),
    .Y(_03882_));
 sky130_fd_sc_hd__or2_1 _09976_ (.A(_03860_),
    .B(_03882_),
    .X(_03883_));
 sky130_fd_sc_hd__nand2_1 _09977_ (.A(_03882_),
    .B(_03860_),
    .Y(_03884_));
 sky130_fd_sc_hd__nand2_1 _09978_ (.A(_03883_),
    .B(_03884_),
    .Y(_03885_));
 sky130_fd_sc_hd__nand3_2 _09979_ (.A(_03859_),
    .B(_02785_),
    .C(_03050_),
    .Y(_03886_));
 sky130_fd_sc_hd__nand2_1 _09980_ (.A(_02619_),
    .B(_03876_),
    .Y(_03887_));
 sky130_fd_sc_hd__or2_1 _09981_ (.A(_03880_),
    .B(_03887_),
    .X(_03888_));
 sky130_fd_sc_hd__nand2_1 _09982_ (.A(_02619_),
    .B(_03868_),
    .Y(_03889_));
 sky130_fd_sc_hd__nand2_1 _09983_ (.A(_03877_),
    .B(_03889_),
    .Y(_03890_));
 sky130_fd_sc_hd__nand2_1 _09984_ (.A(_03888_),
    .B(_03890_),
    .Y(_03891_));
 sky130_fd_sc_hd__o21ai_1 _09985_ (.A1(_03886_),
    .A2(_03891_),
    .B1(_03888_),
    .Y(_03892_));
 sky130_fd_sc_hd__inv_2 _09986_ (.A(_03892_),
    .Y(_03893_));
 sky130_fd_sc_hd__nand2_1 _09987_ (.A(_03885_),
    .B(_03893_),
    .Y(_03894_));
 sky130_fd_sc_hd__nand3_1 _09988_ (.A(_03892_),
    .B(_03883_),
    .C(_03884_),
    .Y(_03895_));
 sky130_fd_sc_hd__nand2_1 _09989_ (.A(_03894_),
    .B(_03895_),
    .Y(_03896_));
 sky130_fd_sc_hd__clkbuf_4 _09990_ (.A(_03049_),
    .X(_03897_));
 sky130_fd_sc_hd__inv_2 _09991_ (.A(_03835_),
    .Y(_03898_));
 sky130_fd_sc_hd__buf_4 _09992_ (.A(_03898_),
    .X(_03899_));
 sky130_fd_sc_hd__or3_1 _09993_ (.A(_03897_),
    .B(_03205_),
    .C(_03899_),
    .X(_03900_));
 sky130_fd_sc_hd__nand2_1 _09994_ (.A(_03896_),
    .B(_03900_),
    .Y(_03901_));
 sky130_fd_sc_hd__nand3b_1 _09995_ (.A_N(_03900_),
    .B(_03894_),
    .C(_03895_),
    .Y(_03902_));
 sky130_fd_sc_hd__nand2_1 _09996_ (.A(_03901_),
    .B(_03902_),
    .Y(_03903_));
 sky130_fd_sc_hd__or3_1 _09997_ (.A(_02949_),
    .B(_03897_),
    .C(_03899_),
    .X(_03904_));
 sky130_fd_sc_hd__xnor2_1 _09998_ (.A(_03886_),
    .B(_03891_),
    .Y(_03905_));
 sky130_fd_sc_hd__nand3_1 _09999_ (.A(_03835_),
    .B(_02785_),
    .C(_03050_),
    .Y(_03906_));
 sky130_fd_sc_hd__inv_2 _10000_ (.A(_03906_),
    .Y(_03907_));
 sky130_fd_sc_hd__nor2_1 _10001_ (.A(_03049_),
    .B(_02738_),
    .Y(_03908_));
 sky130_fd_sc_hd__nand2_1 _10002_ (.A(_03908_),
    .B(_03859_),
    .Y(_03909_));
 sky130_fd_sc_hd__nand2_1 _10003_ (.A(_03909_),
    .B(_03887_),
    .Y(_03910_));
 sky130_fd_sc_hd__nor2_1 _10004_ (.A(_03887_),
    .B(_03909_),
    .Y(_03911_));
 sky130_fd_sc_hd__a21oi_1 _10005_ (.A1(_03907_),
    .A2(_03910_),
    .B1(_03911_),
    .Y(_03912_));
 sky130_fd_sc_hd__nand2_1 _10006_ (.A(_03905_),
    .B(_03912_),
    .Y(_03913_));
 sky130_fd_sc_hd__inv_2 _10007_ (.A(_03913_),
    .Y(_03914_));
 sky130_fd_sc_hd__xor2_1 _10008_ (.A(_03886_),
    .B(_03891_),
    .X(_03915_));
 sky130_fd_sc_hd__inv_2 _10009_ (.A(_03912_),
    .Y(_03916_));
 sky130_fd_sc_hd__nand2_1 _10010_ (.A(_03915_),
    .B(_03916_),
    .Y(_03917_));
 sky130_fd_sc_hd__o21a_1 _10011_ (.A1(_03904_),
    .A2(_03914_),
    .B1(_03917_),
    .X(_03918_));
 sky130_fd_sc_hd__nor2_1 _10012_ (.A(_03903_),
    .B(_03918_),
    .Y(_03919_));
 sky130_fd_sc_hd__nand2_1 _10013_ (.A(_03918_),
    .B(_03903_),
    .Y(_03920_));
 sky130_fd_sc_hd__inv_2 _10014_ (.A(_03920_),
    .Y(_03921_));
 sky130_fd_sc_hd__nor2_1 _10015_ (.A(_03919_),
    .B(_03921_),
    .Y(_03922_));
 sky130_fd_sc_hd__nand2_1 _10016_ (.A(_03902_),
    .B(_03895_),
    .Y(_03923_));
 sky130_fd_sc_hd__inv_2 _10017_ (.A(_03923_),
    .Y(_03924_));
 sky130_fd_sc_hd__or3_1 _10018_ (.A(_03897_),
    .B(_03350_),
    .C(_03898_),
    .X(_03925_));
 sky130_fd_sc_hd__nand2_1 _10019_ (.A(_03883_),
    .B(_03878_),
    .Y(_03926_));
 sky130_fd_sc_hd__nand3_1 _10020_ (.A(_03858_),
    .B(_03050_),
    .C(_03020_),
    .Y(_03927_));
 sky130_fd_sc_hd__nand2_1 _10021_ (.A(_02963_),
    .B(_03868_),
    .Y(_03928_));
 sky130_fd_sc_hd__or2_1 _10022_ (.A(_03879_),
    .B(_03928_),
    .X(_03929_));
 sky130_fd_sc_hd__nand2_1 _10023_ (.A(_02963_),
    .B(_03876_),
    .Y(_03930_));
 sky130_fd_sc_hd__nand2_1 _10024_ (.A(_03930_),
    .B(_03869_),
    .Y(_03931_));
 sky130_fd_sc_hd__nand2_1 _10025_ (.A(_03929_),
    .B(_03931_),
    .Y(_03932_));
 sky130_fd_sc_hd__or2_1 _10026_ (.A(_03927_),
    .B(_03932_),
    .X(_03933_));
 sky130_fd_sc_hd__nand2_1 _10027_ (.A(_03932_),
    .B(_03927_),
    .Y(_03934_));
 sky130_fd_sc_hd__nand3_1 _10028_ (.A(_03926_),
    .B(_03933_),
    .C(_03934_),
    .Y(_03935_));
 sky130_fd_sc_hd__nand2_1 _10029_ (.A(_03933_),
    .B(_03934_),
    .Y(_03936_));
 sky130_fd_sc_hd__nand3_1 _10030_ (.A(_03936_),
    .B(_03878_),
    .C(_03883_),
    .Y(_03937_));
 sky130_fd_sc_hd__nand3b_1 _10031_ (.A_N(_03925_),
    .B(_03935_),
    .C(_03937_),
    .Y(_03938_));
 sky130_fd_sc_hd__nand2_1 _10032_ (.A(_03937_),
    .B(_03935_),
    .Y(_03939_));
 sky130_fd_sc_hd__nand2_1 _10033_ (.A(_03939_),
    .B(_03925_),
    .Y(_03940_));
 sky130_fd_sc_hd__nand3_1 _10034_ (.A(_03924_),
    .B(_03938_),
    .C(_03940_),
    .Y(_03941_));
 sky130_fd_sc_hd__nand2_1 _10035_ (.A(_03940_),
    .B(_03938_),
    .Y(_03942_));
 sky130_fd_sc_hd__nand2_1 _10036_ (.A(_03942_),
    .B(_03923_),
    .Y(_03943_));
 sky130_fd_sc_hd__nand2_1 _10037_ (.A(_03941_),
    .B(_03943_),
    .Y(_03944_));
 sky130_fd_sc_hd__inv_2 _10038_ (.A(_03910_),
    .Y(_03945_));
 sky130_fd_sc_hd__nor2_1 _10039_ (.A(_03911_),
    .B(_03945_),
    .Y(_03946_));
 sky130_fd_sc_hd__xor2_1 _10040_ (.A(_03906_),
    .B(_03946_),
    .X(_03947_));
 sky130_fd_sc_hd__inv_2 _10041_ (.A(_03947_),
    .Y(_03948_));
 sky130_fd_sc_hd__or3b_1 _10042_ (.A(_03897_),
    .B(_03899_),
    .C_N(_02620_),
    .X(_03949_));
 sky130_fd_sc_hd__nor2_1 _10043_ (.A(_03909_),
    .B(_03949_),
    .Y(_03950_));
 sky130_fd_sc_hd__nand2_1 _10044_ (.A(_03948_),
    .B(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__nand2_1 _10045_ (.A(_03917_),
    .B(_03913_),
    .Y(_03952_));
 sky130_fd_sc_hd__nand2_1 _10046_ (.A(_03952_),
    .B(_03904_),
    .Y(_03953_));
 sky130_fd_sc_hd__nand3b_1 _10047_ (.A_N(_03904_),
    .B(_03917_),
    .C(_03913_),
    .Y(_03954_));
 sky130_fd_sc_hd__nand2_1 _10048_ (.A(_03953_),
    .B(_03954_),
    .Y(_03955_));
 sky130_fd_sc_hd__nor2_2 _10049_ (.A(_03951_),
    .B(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__nand3_1 _10050_ (.A(_03922_),
    .B(_03944_),
    .C(_03956_),
    .Y(_03957_));
 sky130_fd_sc_hd__nand2_1 _10051_ (.A(_03942_),
    .B(_03924_),
    .Y(_03958_));
 sky130_fd_sc_hd__nor2_1 _10052_ (.A(_03924_),
    .B(_03942_),
    .Y(_03959_));
 sky130_fd_sc_hd__a21oi_1 _10053_ (.A1(_03958_),
    .A2(_03919_),
    .B1(_03959_),
    .Y(_03960_));
 sky130_fd_sc_hd__nand2_1 _10054_ (.A(_03957_),
    .B(_03960_),
    .Y(_03961_));
 sky130_fd_sc_hd__nand3_1 _10055_ (.A(_03858_),
    .B(_03050_),
    .C(_03421_),
    .Y(_03962_));
 sky130_fd_sc_hd__nand2_1 _10056_ (.A(_03019_),
    .B(_03868_),
    .Y(_03963_));
 sky130_fd_sc_hd__or2_1 _10057_ (.A(_03930_),
    .B(_03963_),
    .X(_03964_));
 sky130_fd_sc_hd__nand2_1 _10058_ (.A(_03019_),
    .B(_03876_),
    .Y(_03965_));
 sky130_fd_sc_hd__nand2_1 _10059_ (.A(_03965_),
    .B(_03928_),
    .Y(_03966_));
 sky130_fd_sc_hd__nand2_1 _10060_ (.A(_03964_),
    .B(_03966_),
    .Y(_03967_));
 sky130_fd_sc_hd__or2_1 _10061_ (.A(_03962_),
    .B(_03967_),
    .X(_03968_));
 sky130_fd_sc_hd__nand2_1 _10062_ (.A(_03967_),
    .B(_03962_),
    .Y(_03969_));
 sky130_fd_sc_hd__nand2_1 _10063_ (.A(_03968_),
    .B(_03969_),
    .Y(_03970_));
 sky130_fd_sc_hd__and2_1 _10064_ (.A(_03933_),
    .B(_03929_),
    .X(_03971_));
 sky130_fd_sc_hd__or2_1 _10065_ (.A(_03970_),
    .B(_03971_),
    .X(_03972_));
 sky130_fd_sc_hd__nand2_1 _10066_ (.A(_03971_),
    .B(_03970_),
    .Y(_03973_));
 sky130_fd_sc_hd__nand2_1 _10067_ (.A(_03972_),
    .B(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__or3_1 _10068_ (.A(_03049_),
    .B(_03507_),
    .C(_03898_),
    .X(_03975_));
 sky130_fd_sc_hd__nand2_1 _10069_ (.A(_03974_),
    .B(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hd__inv_2 _10070_ (.A(_03975_),
    .Y(_03977_));
 sky130_fd_sc_hd__nand3_1 _10071_ (.A(_03972_),
    .B(_03973_),
    .C(_03977_),
    .Y(_03978_));
 sky130_fd_sc_hd__nand2_1 _10072_ (.A(_03976_),
    .B(_03978_),
    .Y(_03979_));
 sky130_fd_sc_hd__nand2_1 _10073_ (.A(_03938_),
    .B(_03935_),
    .Y(_03980_));
 sky130_fd_sc_hd__inv_2 _10074_ (.A(_03980_),
    .Y(_03981_));
 sky130_fd_sc_hd__nand2_1 _10075_ (.A(_03979_),
    .B(_03981_),
    .Y(_03982_));
 sky130_fd_sc_hd__nand3_2 _10076_ (.A(_03976_),
    .B(_03978_),
    .C(_03980_),
    .Y(_03983_));
 sky130_fd_sc_hd__nand2_1 _10077_ (.A(_03982_),
    .B(_03983_),
    .Y(_03984_));
 sky130_fd_sc_hd__inv_2 _10078_ (.A(_03984_),
    .Y(_03985_));
 sky130_fd_sc_hd__nand2_1 _10079_ (.A(_03961_),
    .B(_03985_),
    .Y(_03986_));
 sky130_fd_sc_hd__nand2_1 _10080_ (.A(_03986_),
    .B(_03983_),
    .Y(_03987_));
 sky130_fd_sc_hd__nand3_1 _10081_ (.A(_03858_),
    .B(_03506_),
    .C(_03050_),
    .Y(_03988_));
 sky130_fd_sc_hd__nand2_1 _10082_ (.A(_03349_),
    .B(_03868_),
    .Y(_03989_));
 sky130_fd_sc_hd__or2_1 _10083_ (.A(_03965_),
    .B(_03989_),
    .X(_03990_));
 sky130_fd_sc_hd__nand2_1 _10084_ (.A(_03421_),
    .B(_03876_),
    .Y(_03991_));
 sky130_fd_sc_hd__nand2_1 _10085_ (.A(_03991_),
    .B(_03963_),
    .Y(_03992_));
 sky130_fd_sc_hd__nand2_1 _10086_ (.A(_03990_),
    .B(_03992_),
    .Y(_03993_));
 sky130_fd_sc_hd__or2_1 _10087_ (.A(_03988_),
    .B(_03993_),
    .X(_03994_));
 sky130_fd_sc_hd__nand2_1 _10088_ (.A(_03993_),
    .B(_03988_),
    .Y(_03995_));
 sky130_fd_sc_hd__nand2_1 _10089_ (.A(_03994_),
    .B(_03995_),
    .Y(_03996_));
 sky130_fd_sc_hd__a21o_1 _10090_ (.A1(_03964_),
    .A2(_03968_),
    .B1(_03996_),
    .X(_03997_));
 sky130_fd_sc_hd__nand3_1 _10091_ (.A(_03996_),
    .B(_03964_),
    .C(_03968_),
    .Y(_03998_));
 sky130_fd_sc_hd__nand2_1 _10092_ (.A(_03997_),
    .B(_03998_),
    .Y(_03999_));
 sky130_fd_sc_hd__or3_1 _10093_ (.A(_03897_),
    .B(_03899_),
    .C(_03685_),
    .X(_04000_));
 sky130_fd_sc_hd__nand2_1 _10094_ (.A(_03999_),
    .B(_04000_),
    .Y(_04001_));
 sky130_fd_sc_hd__nand3b_2 _10095_ (.A_N(_04000_),
    .B(_03997_),
    .C(_03998_),
    .Y(_04002_));
 sky130_fd_sc_hd__nand2_1 _10096_ (.A(_04001_),
    .B(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__nand2_1 _10097_ (.A(_03978_),
    .B(_03972_),
    .Y(_04004_));
 sky130_fd_sc_hd__inv_2 _10098_ (.A(_04004_),
    .Y(_04005_));
 sky130_fd_sc_hd__nand2_1 _10099_ (.A(_04003_),
    .B(_04005_),
    .Y(_04006_));
 sky130_fd_sc_hd__nand3_2 _10100_ (.A(_04004_),
    .B(_04001_),
    .C(_04002_),
    .Y(_04007_));
 sky130_fd_sc_hd__nand2_1 _10101_ (.A(_04006_),
    .B(_04007_),
    .Y(_04008_));
 sky130_fd_sc_hd__inv_2 _10102_ (.A(_04008_),
    .Y(_04009_));
 sky130_fd_sc_hd__nand2_1 _10103_ (.A(_03987_),
    .B(_04009_),
    .Y(_04010_));
 sky130_fd_sc_hd__and2_1 _10104_ (.A(_04002_),
    .B(_03997_),
    .X(_04011_));
 sky130_fd_sc_hd__and2_1 _10105_ (.A(_03994_),
    .B(_03990_),
    .X(_04012_));
 sky130_fd_sc_hd__nand2_1 _10106_ (.A(_03505_),
    .B(_03876_),
    .Y(_04013_));
 sky130_fd_sc_hd__or2_1 _10107_ (.A(_03989_),
    .B(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__nand2_1 _10108_ (.A(_04013_),
    .B(_03989_),
    .Y(_04015_));
 sky130_fd_sc_hd__nand2_1 _10109_ (.A(_04014_),
    .B(_04015_),
    .Y(_04016_));
 sky130_fd_sc_hd__nand3_1 _10110_ (.A(_03652_),
    .B(_03745_),
    .C(_03859_),
    .Y(_04017_));
 sky130_fd_sc_hd__or2_1 _10111_ (.A(_04016_),
    .B(_04017_),
    .X(_04018_));
 sky130_fd_sc_hd__nand2_1 _10112_ (.A(_04017_),
    .B(_04016_),
    .Y(_04019_));
 sky130_fd_sc_hd__nand2_1 _10113_ (.A(_04018_),
    .B(_04019_),
    .Y(_04020_));
 sky130_fd_sc_hd__or2_1 _10114_ (.A(_04012_),
    .B(_04020_),
    .X(_04021_));
 sky130_fd_sc_hd__nand2_1 _10115_ (.A(_04020_),
    .B(_04012_),
    .Y(_04022_));
 sky130_fd_sc_hd__nand2_1 _10116_ (.A(_04021_),
    .B(_04022_),
    .Y(_04023_));
 sky130_fd_sc_hd__nand3b_1 _10117_ (.A_N(_04023_),
    .B(_03790_),
    .C(_03835_),
    .Y(_04024_));
 sky130_fd_sc_hd__inv_2 _10118_ (.A(_03789_),
    .Y(_04025_));
 sky130_fd_sc_hd__o21ai_1 _10119_ (.A1(_04025_),
    .A2(_03899_),
    .B1(_04023_),
    .Y(_04026_));
 sky130_fd_sc_hd__nand2_1 _10120_ (.A(_04024_),
    .B(_04026_),
    .Y(_04027_));
 sky130_fd_sc_hd__or2_1 _10121_ (.A(_04011_),
    .B(_04027_),
    .X(_04028_));
 sky130_fd_sc_hd__nand2_1 _10122_ (.A(_04027_),
    .B(_04011_),
    .Y(_04029_));
 sky130_fd_sc_hd__nand2_1 _10123_ (.A(_04028_),
    .B(_04029_),
    .Y(_04030_));
 sky130_fd_sc_hd__nand3_1 _10124_ (.A(_04010_),
    .B(_04007_),
    .C(_04030_),
    .Y(_04031_));
 sky130_fd_sc_hd__nor2_1 _10125_ (.A(_03984_),
    .B(_04008_),
    .Y(_04032_));
 sky130_fd_sc_hd__and2_1 _10126_ (.A(_03922_),
    .B(_03944_),
    .X(_04033_));
 sky130_fd_sc_hd__nand3_1 _10127_ (.A(_04032_),
    .B(_03956_),
    .C(_04033_),
    .Y(_04034_));
 sky130_fd_sc_hd__nand3b_1 _10128_ (.A_N(_03960_),
    .B(_04009_),
    .C(_03985_),
    .Y(_04035_));
 sky130_fd_sc_hd__inv_2 _10129_ (.A(_04006_),
    .Y(_04036_));
 sky130_fd_sc_hd__o21a_1 _10130_ (.A1(_03983_),
    .A2(_04036_),
    .B1(_04007_),
    .X(_04037_));
 sky130_fd_sc_hd__nand3_1 _10131_ (.A(_04034_),
    .B(_04035_),
    .C(_04037_),
    .Y(_04038_));
 sky130_fd_sc_hd__inv_2 _10132_ (.A(_04030_),
    .Y(_04039_));
 sky130_fd_sc_hd__nand2_2 _10133_ (.A(_04038_),
    .B(_04039_),
    .Y(_04040_));
 sky130_fd_sc_hd__nand2_1 _10134_ (.A(_04031_),
    .B(_04040_),
    .Y(_04041_));
 sky130_fd_sc_hd__buf_4 _10135_ (.A(_02560_),
    .X(_04042_));
 sky130_fd_sc_hd__mux2_1 _10136_ (.A0(\H[0][13] ),
    .A1(\H[1][13] ),
    .S(_02545_),
    .X(_04043_));
 sky130_fd_sc_hd__nand2_1 _10137_ (.A(_03152_),
    .B(\H[2][13] ),
    .Y(_04044_));
 sky130_fd_sc_hd__buf_4 _10138_ (.A(_03135_),
    .X(_04045_));
 sky130_fd_sc_hd__a21oi_1 _10139_ (.A1(_02567_),
    .A2(\H[3][13] ),
    .B1(_04045_),
    .Y(_04046_));
 sky130_fd_sc_hd__a2bb2o_2 _10140_ (.A1_N(_04042_),
    .A2_N(_04043_),
    .B1(_04044_),
    .B2(_04046_),
    .X(_04047_));
 sky130_fd_sc_hd__or2_2 _10141_ (.A(_00588_),
    .B(_04047_),
    .X(_04048_));
 sky130_fd_sc_hd__nor2_2 _10142_ (.A(_03758_),
    .B(_04048_),
    .Y(_04049_));
 sky130_fd_sc_hd__inv_2 _10143_ (.A(_04049_),
    .Y(_04050_));
 sky130_fd_sc_hd__nor2_1 _10144_ (.A(_03115_),
    .B(_04050_),
    .Y(_04051_));
 sky130_fd_sc_hd__inv_2 _10145_ (.A(_04051_),
    .Y(_04052_));
 sky130_fd_sc_hd__inv_2 _10146_ (.A(\Qset[1][14] ),
    .Y(_04053_));
 sky130_fd_sc_hd__a21oi_1 _10147_ (.A1(_03136_),
    .A2(\Qset[0][14] ),
    .B1(_02526_),
    .Y(_04054_));
 sky130_fd_sc_hd__o21ai_1 _10148_ (.A1(_03152_),
    .A2(_04053_),
    .B1(_04054_),
    .Y(_04055_));
 sky130_fd_sc_hd__a21oi_1 _10149_ (.A1(_03157_),
    .A2(\Qset[3][14] ),
    .B1(_02535_),
    .Y(_04056_));
 sky130_fd_sc_hd__o21ai_1 _10150_ (.A1(_02565_),
    .A2(_02476_),
    .B1(_04056_),
    .Y(_04057_));
 sky130_fd_sc_hd__nand2_2 _10151_ (.A(_04055_),
    .B(_04057_),
    .Y(_04058_));
 sky130_fd_sc_hd__o21ai_1 _10152_ (.A1(_02162_),
    .A2(_04058_),
    .B1(_02796_),
    .Y(_04059_));
 sky130_fd_sc_hd__nand2_1 _10153_ (.A(_02523_),
    .B(_02483_),
    .Y(_04060_));
 sky130_fd_sc_hd__o211a_1 _10154_ (.A1(\Oset[3][14] ),
    .A2(_02787_),
    .B1(_02525_),
    .C1(_04060_),
    .X(_04061_));
 sky130_fd_sc_hd__nand2_1 _10155_ (.A(_02523_),
    .B(_02486_),
    .Y(_04062_));
 sky130_fd_sc_hd__o211a_1 _10156_ (.A1(\Oset[1][14] ),
    .A2(_02523_),
    .B1(_02535_),
    .C1(_04062_),
    .X(_04063_));
 sky130_fd_sc_hd__nor2_2 _10157_ (.A(_04061_),
    .B(_04063_),
    .Y(_04064_));
 sky130_fd_sc_hd__nand2_1 _10158_ (.A(_04064_),
    .B(_02552_),
    .Y(_04065_));
 sky130_fd_sc_hd__a31o_1 _10159_ (.A1(_04059_),
    .A2(_04065_),
    .A3(_01155_),
    .B1(_03095_),
    .X(_04066_));
 sky130_fd_sc_hd__nor2_1 _10160_ (.A(_02565_),
    .B(\H[0][14] ),
    .Y(_04067_));
 sky130_fd_sc_hd__nor2_1 _10161_ (.A(\H[1][14] ),
    .B(_03152_),
    .Y(_04068_));
 sky130_fd_sc_hd__nor2_1 _10162_ (.A(_03157_),
    .B(\H[2][14] ),
    .Y(_04069_));
 sky130_fd_sc_hd__a211o_1 _10163_ (.A1(_02490_),
    .A2(_03157_),
    .B1(_03135_),
    .C1(_04069_),
    .X(_04070_));
 sky130_fd_sc_hd__o31a_2 _10164_ (.A1(_02560_),
    .A2(_04067_),
    .A3(_04068_),
    .B1(_04070_),
    .X(_04071_));
 sky130_fd_sc_hd__a21oi_1 _10165_ (.A1(_04071_),
    .A2(_02573_),
    .B1(_00588_),
    .Y(_04072_));
 sky130_fd_sc_hd__nand2_4 _10166_ (.A(_04066_),
    .B(_04072_),
    .Y(_04073_));
 sky130_fd_sc_hd__nor2_4 _10167_ (.A(_02556_),
    .B(_04073_),
    .Y(_04074_));
 sky130_fd_sc_hd__nand2_1 _10168_ (.A(_04074_),
    .B(_02620_),
    .Y(_04075_));
 sky130_fd_sc_hd__inv_2 _10169_ (.A(\Qset[1][15] ),
    .Y(_04076_));
 sky130_fd_sc_hd__a21oi_1 _10170_ (.A1(_03136_),
    .A2(\Qset[0][15] ),
    .B1(_02526_),
    .Y(_04077_));
 sky130_fd_sc_hd__o21ai_2 _10171_ (.A1(_03136_),
    .A2(_04076_),
    .B1(_04077_),
    .Y(_04078_));
 sky130_fd_sc_hd__a21oi_1 _10172_ (.A1(_03157_),
    .A2(\Qset[3][15] ),
    .B1(_02535_),
    .Y(_04079_));
 sky130_fd_sc_hd__o21ai_2 _10173_ (.A1(_02565_),
    .A2(_02500_),
    .B1(_04079_),
    .Y(_04080_));
 sky130_fd_sc_hd__a31o_1 _10174_ (.A1(_04078_),
    .A2(_04080_),
    .A3(_00581_),
    .B1(_02871_),
    .X(_04081_));
 sky130_fd_sc_hd__a21oi_1 _10175_ (.A1(_02529_),
    .A2(\Oset[3][15] ),
    .B1(_02535_),
    .Y(_04082_));
 sky130_fd_sc_hd__nand2_1 _10176_ (.A(_02523_),
    .B(\Oset[2][15] ),
    .Y(_04083_));
 sky130_fd_sc_hd__a21oi_1 _10177_ (.A1(_02523_),
    .A2(\Oset[0][15] ),
    .B1(_02525_),
    .Y(_04084_));
 sky130_fd_sc_hd__nand2_1 _10178_ (.A(_02545_),
    .B(\Oset[1][15] ),
    .Y(_04085_));
 sky130_fd_sc_hd__a22o_2 _10179_ (.A1(_04082_),
    .A2(_04083_),
    .B1(_04084_),
    .B2(_04085_),
    .X(_04086_));
 sky130_fd_sc_hd__nand2_1 _10180_ (.A(_04086_),
    .B(_02552_),
    .Y(_04087_));
 sky130_fd_sc_hd__a31o_1 _10181_ (.A1(_04081_),
    .A2(_01155_),
    .A3(_04087_),
    .B1(_03066_),
    .X(_04088_));
 sky130_fd_sc_hd__nand2_1 _10182_ (.A(_03152_),
    .B(_02514_),
    .Y(_04089_));
 sky130_fd_sc_hd__o211a_1 _10183_ (.A1(\H[1][15] ),
    .A2(_03152_),
    .B1(_03135_),
    .C1(_04089_),
    .X(_04090_));
 sky130_fd_sc_hd__or2_1 _10184_ (.A(_02529_),
    .B(\H[2][15] ),
    .X(_04091_));
 sky130_fd_sc_hd__o211a_1 _10185_ (.A1(_03152_),
    .A2(\H[3][15] ),
    .B1(_02560_),
    .C1(_04091_),
    .X(_04092_));
 sky130_fd_sc_hd__nor2_2 _10186_ (.A(_04090_),
    .B(_04092_),
    .Y(_04093_));
 sky130_fd_sc_hd__a21oi_1 _10187_ (.A1(_04093_),
    .A2(_02573_),
    .B1(_00588_),
    .Y(_04094_));
 sky130_fd_sc_hd__nand2_4 _10188_ (.A(_04088_),
    .B(_04094_),
    .Y(_04095_));
 sky130_fd_sc_hd__nor2_4 _10189_ (.A(_02556_),
    .B(_04095_),
    .Y(_04096_));
 sky130_fd_sc_hd__nand2_1 _10190_ (.A(_04096_),
    .B(_02687_),
    .Y(_04097_));
 sky130_fd_sc_hd__a22o_1 _10191_ (.A1(_04074_),
    .A2(_02687_),
    .B1(_04096_),
    .B2(_02620_),
    .X(_04098_));
 sky130_fd_sc_hd__o21ai_1 _10192_ (.A1(_04075_),
    .A2(_04097_),
    .B1(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__or2_1 _10193_ (.A(_04052_),
    .B(_04099_),
    .X(_04100_));
 sky130_fd_sc_hd__nand2_1 _10194_ (.A(_04099_),
    .B(_04052_),
    .Y(_04101_));
 sky130_fd_sc_hd__nand2_1 _10195_ (.A(_04100_),
    .B(_04101_),
    .Y(_04102_));
 sky130_fd_sc_hd__mux2_1 _10196_ (.A0(\H[0][12] ),
    .A1(\H[1][12] ),
    .S(_02567_),
    .X(_04103_));
 sky130_fd_sc_hd__nand2_1 _10197_ (.A(_03152_),
    .B(\H[2][12] ),
    .Y(_04104_));
 sky130_fd_sc_hd__buf_6 _10198_ (.A(_02567_),
    .X(_04105_));
 sky130_fd_sc_hd__a21oi_1 _10199_ (.A1(_04105_),
    .A2(\H[3][12] ),
    .B1(_04045_),
    .Y(_04106_));
 sky130_fd_sc_hd__a2bb2o_1 _10200_ (.A1_N(_04042_),
    .A2_N(_04103_),
    .B1(_04104_),
    .B2(_04106_),
    .X(_04107_));
 sky130_fd_sc_hd__or2_2 _10201_ (.A(_00589_),
    .B(_04107_),
    .X(_04108_));
 sky130_fd_sc_hd__nor2_2 _10202_ (.A(_03758_),
    .B(_04108_),
    .Y(_04109_));
 sky130_fd_sc_hd__inv_2 _10203_ (.A(_04109_),
    .Y(_04110_));
 sky130_fd_sc_hd__nor2_1 _10204_ (.A(_03115_),
    .B(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__nand2_1 _10205_ (.A(_04049_),
    .B(_02687_),
    .Y(_04112_));
 sky130_fd_sc_hd__nand2_1 _10206_ (.A(_04075_),
    .B(_04112_),
    .Y(_04113_));
 sky130_fd_sc_hd__nand2_1 _10207_ (.A(_04049_),
    .B(_02620_),
    .Y(_04114_));
 sky130_fd_sc_hd__nand2_1 _10208_ (.A(_04074_),
    .B(_02687_),
    .Y(_04115_));
 sky130_fd_sc_hd__o2bb2a_1 _10209_ (.A1_N(_04111_),
    .A2_N(_04113_),
    .B1(_04114_),
    .B2(_04115_),
    .X(_04116_));
 sky130_fd_sc_hd__nand2_1 _10210_ (.A(_04102_),
    .B(_04116_),
    .Y(_04117_));
 sky130_fd_sc_hd__nor2_1 _10211_ (.A(_02949_),
    .B(_04110_),
    .Y(_04118_));
 sky130_fd_sc_hd__nand3b_1 _10212_ (.A_N(_04116_),
    .B(_04100_),
    .C(_04101_),
    .Y(_04119_));
 sky130_fd_sc_hd__a21boi_1 _10213_ (.A1(_04117_),
    .A2(_04118_),
    .B1_N(_04119_),
    .Y(_04120_));
 sky130_fd_sc_hd__nor2_1 _10214_ (.A(_04075_),
    .B(_04097_),
    .Y(_04121_));
 sky130_fd_sc_hd__a21oi_1 _10215_ (.A1(_04098_),
    .A2(_04051_),
    .B1(_04121_),
    .Y(_04122_));
 sky130_fd_sc_hd__nor2_1 _10216_ (.A(_02949_),
    .B(_04050_),
    .Y(_04123_));
 sky130_fd_sc_hd__nand2_1 _10217_ (.A(_04096_),
    .B(_02785_),
    .Y(_04124_));
 sky130_fd_sc_hd__nand2_1 _10218_ (.A(_04074_),
    .B(_02785_),
    .Y(_04125_));
 sky130_fd_sc_hd__nand2_1 _10219_ (.A(_04097_),
    .B(_04125_),
    .Y(_04126_));
 sky130_fd_sc_hd__o21a_1 _10220_ (.A1(_04115_),
    .A2(_04124_),
    .B1(_04126_),
    .X(_04127_));
 sky130_fd_sc_hd__or2_1 _10221_ (.A(_04123_),
    .B(_04127_),
    .X(_04128_));
 sky130_fd_sc_hd__nand2_1 _10222_ (.A(_04127_),
    .B(_04123_),
    .Y(_04129_));
 sky130_fd_sc_hd__nand2_1 _10223_ (.A(_04128_),
    .B(_04129_),
    .Y(_04130_));
 sky130_fd_sc_hd__nor2_1 _10224_ (.A(_04122_),
    .B(_04130_),
    .Y(_04131_));
 sky130_fd_sc_hd__nand2_1 _10225_ (.A(_04130_),
    .B(_04122_),
    .Y(_04132_));
 sky130_fd_sc_hd__inv_2 _10226_ (.A(_04132_),
    .Y(_04133_));
 sky130_fd_sc_hd__nor2_1 _10227_ (.A(_03205_),
    .B(_04110_),
    .Y(_04134_));
 sky130_fd_sc_hd__o21bai_1 _10228_ (.A1(_04131_),
    .A2(_04133_),
    .B1_N(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__nand3b_1 _10229_ (.A_N(_04131_),
    .B(_04134_),
    .C(_04132_),
    .Y(_04136_));
 sky130_fd_sc_hd__nand2_1 _10230_ (.A(_04135_),
    .B(_04136_),
    .Y(_04137_));
 sky130_fd_sc_hd__nor2_1 _10231_ (.A(_04120_),
    .B(_04137_),
    .Y(_04138_));
 sky130_fd_sc_hd__nand2_1 _10232_ (.A(_04137_),
    .B(_04120_),
    .Y(_04139_));
 sky130_fd_sc_hd__inv_2 _10233_ (.A(_04139_),
    .Y(_04140_));
 sky130_fd_sc_hd__nand2_1 _10234_ (.A(_04117_),
    .B(_04119_),
    .Y(_04141_));
 sky130_fd_sc_hd__o21ai_1 _10235_ (.A1(_02949_),
    .A2(_04110_),
    .B1(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__nand3_1 _10236_ (.A(_04117_),
    .B(_04119_),
    .C(_04118_),
    .Y(_04143_));
 sky130_fd_sc_hd__o21ai_1 _10237_ (.A1(_04114_),
    .A2(_04115_),
    .B1(_04113_),
    .Y(_04144_));
 sky130_fd_sc_hd__xor2_1 _10238_ (.A(_04111_),
    .B(_04144_),
    .X(_04145_));
 sky130_fd_sc_hd__inv_2 _10239_ (.A(_04145_),
    .Y(_04146_));
 sky130_fd_sc_hd__nand2_2 _10240_ (.A(_04109_),
    .B(_02620_),
    .Y(_04147_));
 sky130_fd_sc_hd__nor2_1 _10241_ (.A(_04112_),
    .B(_04147_),
    .Y(_04148_));
 sky130_fd_sc_hd__nand2_1 _10242_ (.A(_04146_),
    .B(_04148_),
    .Y(_04149_));
 sky130_fd_sc_hd__inv_2 _10243_ (.A(_04149_),
    .Y(_04150_));
 sky130_fd_sc_hd__nand3_2 _10244_ (.A(_04142_),
    .B(_04143_),
    .C(_04150_),
    .Y(_04151_));
 sky130_fd_sc_hd__o21ai_1 _10245_ (.A1(_04138_),
    .A2(_04140_),
    .B1(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__inv_2 _10246_ (.A(_04151_),
    .Y(_04153_));
 sky130_fd_sc_hd__nand3b_1 _10247_ (.A_N(_04138_),
    .B(_04153_),
    .C(_04139_),
    .Y(_04154_));
 sky130_fd_sc_hd__nand2_1 _10248_ (.A(_04152_),
    .B(_04154_),
    .Y(_04155_));
 sky130_fd_sc_hd__nand2_1 _10249_ (.A(_04041_),
    .B(_04155_),
    .Y(_04156_));
 sky130_fd_sc_hd__nand3b_2 _10250_ (.A_N(_04155_),
    .B(_04031_),
    .C(_04040_),
    .Y(_04157_));
 sky130_fd_sc_hd__nand2_1 _10251_ (.A(_04156_),
    .B(_04157_),
    .Y(_04158_));
 sky130_fd_sc_hd__inv_2 _10252_ (.A(_04158_),
    .Y(_04159_));
 sky130_fd_sc_hd__nand3_1 _10253_ (.A(_03957_),
    .B(_03984_),
    .C(_03960_),
    .Y(_04160_));
 sky130_fd_sc_hd__or2_1 _10254_ (.A(_04148_),
    .B(_04146_),
    .X(_04161_));
 sky130_fd_sc_hd__nand2_1 _10255_ (.A(_04161_),
    .B(_04149_),
    .Y(_04162_));
 sky130_fd_sc_hd__a21boi_1 _10256_ (.A1(_03986_),
    .A2(_04160_),
    .B1_N(_04162_),
    .Y(_04163_));
 sky130_fd_sc_hd__a21oi_1 _10257_ (.A1(_03920_),
    .A2(_03956_),
    .B1(_03919_),
    .Y(_04164_));
 sky130_fd_sc_hd__inv_2 _10258_ (.A(_04164_),
    .Y(_04165_));
 sky130_fd_sc_hd__nand2_1 _10259_ (.A(_04165_),
    .B(_03944_),
    .Y(_04166_));
 sky130_fd_sc_hd__and2_1 _10260_ (.A(_03942_),
    .B(_03924_),
    .X(_04167_));
 sky130_fd_sc_hd__o21ai_1 _10261_ (.A1(_03959_),
    .A2(_04167_),
    .B1(_04164_),
    .Y(_04168_));
 sky130_fd_sc_hd__nand2_1 _10262_ (.A(_04166_),
    .B(_04168_),
    .Y(_04169_));
 sky130_fd_sc_hd__o21ai_1 _10263_ (.A1(_02738_),
    .A2(_04110_),
    .B1(_04114_),
    .Y(_04170_));
 sky130_fd_sc_hd__o21ai_1 _10264_ (.A1(_04112_),
    .A2(_04147_),
    .B1(_04170_),
    .Y(_04171_));
 sky130_fd_sc_hd__nand2_1 _10265_ (.A(_04169_),
    .B(_04171_),
    .Y(_04172_));
 sky130_fd_sc_hd__o21bai_1 _10266_ (.A1(_03919_),
    .A2(_03921_),
    .B1_N(_03956_),
    .Y(_04173_));
 sky130_fd_sc_hd__nand2_1 _10267_ (.A(_03922_),
    .B(_03956_),
    .Y(_04174_));
 sky130_fd_sc_hd__nand2_1 _10268_ (.A(_04173_),
    .B(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__nor2_1 _10269_ (.A(_04147_),
    .B(_04175_),
    .Y(_04176_));
 sky130_fd_sc_hd__nor2_1 _10270_ (.A(_04171_),
    .B(_04169_),
    .Y(_04177_));
 sky130_fd_sc_hd__a21oi_1 _10271_ (.A1(_04172_),
    .A2(_04176_),
    .B1(_04177_),
    .Y(_04178_));
 sky130_fd_sc_hd__nand2_1 _10272_ (.A(_03986_),
    .B(_04160_),
    .Y(_04179_));
 sky130_fd_sc_hd__or2_1 _10273_ (.A(_04162_),
    .B(_04179_),
    .X(_04180_));
 sky130_fd_sc_hd__o21ai_1 _10274_ (.A1(_04163_),
    .A2(_04178_),
    .B1(_04180_),
    .Y(_04181_));
 sky130_fd_sc_hd__nand3_1 _10275_ (.A(_03986_),
    .B(_03983_),
    .C(_04008_),
    .Y(_04182_));
 sky130_fd_sc_hd__nand2_1 _10276_ (.A(_04010_),
    .B(_04182_),
    .Y(_04183_));
 sky130_fd_sc_hd__a21o_1 _10277_ (.A1(_04142_),
    .A2(_04143_),
    .B1(_04150_),
    .X(_04184_));
 sky130_fd_sc_hd__nand2_1 _10278_ (.A(_04184_),
    .B(_04151_),
    .Y(_04185_));
 sky130_fd_sc_hd__inv_2 _10279_ (.A(_04185_),
    .Y(_04186_));
 sky130_fd_sc_hd__nand2_1 _10280_ (.A(_04183_),
    .B(_04186_),
    .Y(_04187_));
 sky130_fd_sc_hd__nand3_1 _10281_ (.A(_04010_),
    .B(_04182_),
    .C(_04185_),
    .Y(_04188_));
 sky130_fd_sc_hd__nand2_1 _10282_ (.A(_04187_),
    .B(_04188_),
    .Y(_04189_));
 sky130_fd_sc_hd__nand2_1 _10283_ (.A(_04181_),
    .B(_04189_),
    .Y(_04190_));
 sky130_fd_sc_hd__or2_1 _10284_ (.A(_04185_),
    .B(_04183_),
    .X(_04191_));
 sky130_fd_sc_hd__nand2_1 _10285_ (.A(_04190_),
    .B(_04191_),
    .Y(_04192_));
 sky130_fd_sc_hd__or2_1 _10286_ (.A(_04159_),
    .B(_04192_),
    .X(_04193_));
 sky130_fd_sc_hd__nand2_1 _10287_ (.A(_04192_),
    .B(_04159_),
    .Y(_04194_));
 sky130_fd_sc_hd__a21o_1 _10288_ (.A1(_04193_),
    .A2(_04194_),
    .B1(_03751_),
    .X(_04195_));
 sky130_fd_sc_hd__buf_4 _10289_ (.A(_03897_),
    .X(_04196_));
 sky130_fd_sc_hd__nand2_1 _10290_ (.A(_04041_),
    .B(_03751_),
    .Y(_04197_));
 sky130_fd_sc_hd__nand3_2 _10291_ (.A(_04195_),
    .B(_04196_),
    .C(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__and2_1 _10292_ (.A(_03655_),
    .B(_03625_),
    .X(_04199_));
 sky130_fd_sc_hd__nand2_1 _10293_ (.A(_03624_),
    .B(_03621_),
    .Y(_04200_));
 sky130_fd_sc_hd__inv_2 _10294_ (.A(_04200_),
    .Y(_04201_));
 sky130_fd_sc_hd__nand2_1 _10295_ (.A(_03506_),
    .B(_03614_),
    .Y(_04202_));
 sky130_fd_sc_hd__nor2_1 _10296_ (.A(_03612_),
    .B(_04202_),
    .Y(_04203_));
 sky130_fd_sc_hd__nand2_1 _10297_ (.A(_03505_),
    .B(_03462_),
    .Y(_04204_));
 sky130_fd_sc_hd__o21ai_1 _10298_ (.A1(_03613_),
    .A2(_03350_),
    .B1(_04204_),
    .Y(_04205_));
 sky130_fd_sc_hd__inv_2 _10299_ (.A(_04205_),
    .Y(_04206_));
 sky130_fd_sc_hd__nor2_1 _10300_ (.A(_04203_),
    .B(_04206_),
    .Y(_04207_));
 sky130_fd_sc_hd__nand2_1 _10301_ (.A(_03651_),
    .B(_03304_),
    .Y(_04208_));
 sky130_fd_sc_hd__inv_2 _10302_ (.A(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__nand2_1 _10303_ (.A(_04207_),
    .B(_04209_),
    .Y(_04210_));
 sky130_fd_sc_hd__o21ai_1 _10304_ (.A1(_04203_),
    .A2(_04206_),
    .B1(_04208_),
    .Y(_04211_));
 sky130_fd_sc_hd__nand2_1 _10305_ (.A(_04210_),
    .B(_04211_),
    .Y(_04212_));
 sky130_fd_sc_hd__or2_1 _10306_ (.A(_04201_),
    .B(_04212_),
    .X(_04213_));
 sky130_fd_sc_hd__nand2_1 _10307_ (.A(_04212_),
    .B(_04201_),
    .Y(_04214_));
 sky130_fd_sc_hd__nand2_1 _10308_ (.A(_04213_),
    .B(_04214_),
    .Y(_04215_));
 sky130_fd_sc_hd__nor2_1 _10309_ (.A(_03897_),
    .B(_02578_),
    .Y(_04216_));
 sky130_fd_sc_hd__nand2_1 _10310_ (.A(_03790_),
    .B(_04216_),
    .Y(_04217_));
 sky130_fd_sc_hd__nand2_1 _10311_ (.A(_04215_),
    .B(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__inv_2 _10312_ (.A(_04217_),
    .Y(_04219_));
 sky130_fd_sc_hd__nand3_1 _10313_ (.A(_04213_),
    .B(_04219_),
    .C(_04214_),
    .Y(_04220_));
 sky130_fd_sc_hd__nand2_1 _10314_ (.A(_04218_),
    .B(_04220_),
    .Y(_04221_));
 sky130_fd_sc_hd__xor2_1 _10315_ (.A(_04199_),
    .B(_04221_),
    .X(_04222_));
 sky130_fd_sc_hd__nand2_1 _10316_ (.A(_03666_),
    .B(_03606_),
    .Y(_04223_));
 sky130_fd_sc_hd__or2_1 _10317_ (.A(_03662_),
    .B(_03659_),
    .X(_04224_));
 sky130_fd_sc_hd__nand2_1 _10318_ (.A(_04223_),
    .B(_04224_),
    .Y(_04225_));
 sky130_fd_sc_hd__nand2_1 _10319_ (.A(_03666_),
    .B(_03518_),
    .Y(_04226_));
 sky130_fd_sc_hd__nor2_1 _10320_ (.A(_04226_),
    .B(_03456_),
    .Y(_04227_));
 sky130_fd_sc_hd__nor2_1 _10321_ (.A(_04225_),
    .B(_04227_),
    .Y(_04228_));
 sky130_fd_sc_hd__nor2_1 _10322_ (.A(_03364_),
    .B(_03266_),
    .Y(_04229_));
 sky130_fd_sc_hd__inv_2 _10323_ (.A(_04226_),
    .Y(_04230_));
 sky130_fd_sc_hd__nand3_1 _10324_ (.A(_04229_),
    .B(_04230_),
    .C(_03270_),
    .Y(_04231_));
 sky130_fd_sc_hd__nand2_1 _10325_ (.A(_04228_),
    .B(_04231_),
    .Y(_04232_));
 sky130_fd_sc_hd__or2_1 _10326_ (.A(_04222_),
    .B(_04232_),
    .X(_04233_));
 sky130_fd_sc_hd__nand2_1 _10327_ (.A(_04232_),
    .B(_04222_),
    .Y(_04234_));
 sky130_fd_sc_hd__nand2_1 _10328_ (.A(_04233_),
    .B(_04234_),
    .Y(_04235_));
 sky130_fd_sc_hd__nand2_1 _10329_ (.A(_03229_),
    .B(_03232_),
    .Y(_04236_));
 sky130_fd_sc_hd__nand2_1 _10330_ (.A(_04235_),
    .B(_04236_),
    .Y(_04237_));
 sky130_fd_sc_hd__inv_2 _10331_ (.A(_04236_),
    .Y(_04238_));
 sky130_fd_sc_hd__nand3_2 _10332_ (.A(_04233_),
    .B(_04238_),
    .C(_04234_),
    .Y(_04239_));
 sky130_fd_sc_hd__and2_1 _10333_ (.A(_04237_),
    .B(_04239_),
    .X(_04240_));
 sky130_fd_sc_hd__nand2_1 _10334_ (.A(_03681_),
    .B(_03674_),
    .Y(_04241_));
 sky130_fd_sc_hd__or2_1 _10335_ (.A(_04240_),
    .B(_04241_),
    .X(_04242_));
 sky130_fd_sc_hd__inv_2 _10336_ (.A(_03949_),
    .Y(_04243_));
 sky130_fd_sc_hd__nand2_1 _10337_ (.A(_04241_),
    .B(_04240_),
    .Y(_04244_));
 sky130_fd_sc_hd__nand3_1 _10338_ (.A(_04242_),
    .B(_04243_),
    .C(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__inv_2 _10339_ (.A(_04245_),
    .Y(_04246_));
 sky130_fd_sc_hd__a21oi_1 _10340_ (.A1(_04242_),
    .A2(_04244_),
    .B1(_04243_),
    .Y(_04247_));
 sky130_fd_sc_hd__or3_2 _10341_ (.A(_04196_),
    .B(_04246_),
    .C(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__nand3_1 _10342_ (.A(_04198_),
    .B(_04248_),
    .C(_00710_),
    .Y(_04249_));
 sky130_fd_sc_hd__o21ai_1 _10343_ (.A1(_00710_),
    .A2(_03835_),
    .B1(_04249_),
    .Y(_04250_));
 sky130_fd_sc_hd__nand2_1 _10344_ (.A(_04250_),
    .B(_02160_),
    .Y(_04251_));
 sky130_fd_sc_hd__o211ai_1 _10345_ (.A1(_00710_),
    .A2(_03835_),
    .B1(_00831_),
    .C1(_04249_),
    .Y(_04252_));
 sky130_fd_sc_hd__nand2_1 _10346_ (.A(_04251_),
    .B(_04252_),
    .Y(_04253_));
 sky130_fd_sc_hd__a21o_1 _10347_ (.A1(_03812_),
    .A2(_03814_),
    .B1(_04253_),
    .X(_04254_));
 sky130_fd_sc_hd__nand3_1 _10348_ (.A(_03812_),
    .B(_03814_),
    .C(_04253_),
    .Y(_04255_));
 sky130_fd_sc_hd__and2_2 _10349_ (.A(_04254_),
    .B(_04255_),
    .X(_04256_));
 sky130_fd_sc_hd__inv_2 _10350_ (.A(_04256_),
    .Y(_04257_));
 sky130_fd_sc_hd__nor2_1 _10351_ (.A(\result_reg_add[8] ),
    .B(_02648_),
    .Y(_04258_));
 sky130_fd_sc_hd__a211o_1 _10352_ (.A1(_04257_),
    .A2(_02649_),
    .B1(_02753_),
    .C1(_04258_),
    .X(_04259_));
 sky130_fd_sc_hd__inv_2 _10353_ (.A(_04259_),
    .Y(_00252_));
 sky130_fd_sc_hd__nand2_1 _10354_ (.A(_04244_),
    .B(_04239_),
    .Y(_04260_));
 sky130_fd_sc_hd__or2_1 _10355_ (.A(_04199_),
    .B(_04221_),
    .X(_04261_));
 sky130_fd_sc_hd__nand2_1 _10356_ (.A(_04234_),
    .B(_04261_),
    .Y(_04262_));
 sky130_fd_sc_hd__a21boi_1 _10357_ (.A1(_04219_),
    .A2(_04214_),
    .B1_N(_04213_),
    .Y(_04263_));
 sky130_fd_sc_hd__inv_2 _10358_ (.A(_04210_),
    .Y(_04264_));
 sky130_fd_sc_hd__nand2_2 _10359_ (.A(_03651_),
    .B(_03614_),
    .Y(_04265_));
 sky130_fd_sc_hd__nor2_1 _10360_ (.A(_04204_),
    .B(_04265_),
    .Y(_04266_));
 sky130_fd_sc_hd__nand2_1 _10361_ (.A(_03651_),
    .B(_03462_),
    .Y(_04267_));
 sky130_fd_sc_hd__nand2_1 _10362_ (.A(_04267_),
    .B(_04202_),
    .Y(_04268_));
 sky130_fd_sc_hd__inv_2 _10363_ (.A(_04268_),
    .Y(_04269_));
 sky130_fd_sc_hd__nor2_2 _10364_ (.A(_03049_),
    .B(_02735_),
    .Y(_04270_));
 sky130_fd_sc_hd__nand2_1 _10365_ (.A(_03789_),
    .B(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__o21ai_1 _10366_ (.A1(_04266_),
    .A2(_04269_),
    .B1(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hd__nor2_1 _10367_ (.A(_04266_),
    .B(_04269_),
    .Y(_04273_));
 sky130_fd_sc_hd__inv_2 _10368_ (.A(_04271_),
    .Y(_04274_));
 sky130_fd_sc_hd__nand2_1 _10369_ (.A(_04273_),
    .B(_04274_),
    .Y(_04275_));
 sky130_fd_sc_hd__nand2_1 _10370_ (.A(_04272_),
    .B(_04275_),
    .Y(_04276_));
 sky130_fd_sc_hd__o21ai_1 _10371_ (.A1(_04203_),
    .A2(_04264_),
    .B1(_04276_),
    .Y(_04277_));
 sky130_fd_sc_hd__nor2_1 _10372_ (.A(_04203_),
    .B(_04264_),
    .Y(_04278_));
 sky130_fd_sc_hd__nand3_1 _10373_ (.A(_04272_),
    .B(_04275_),
    .C(_04278_),
    .Y(_04279_));
 sky130_fd_sc_hd__nand2_1 _10374_ (.A(_04277_),
    .B(_04279_),
    .Y(_04280_));
 sky130_fd_sc_hd__inv_2 _10375_ (.A(_04216_),
    .Y(_04281_));
 sky130_fd_sc_hd__buf_6 _10376_ (.A(_03498_),
    .X(_04282_));
 sky130_fd_sc_hd__buf_6 _10377_ (.A(_04282_),
    .X(_04283_));
 sky130_fd_sc_hd__nor2_1 _10378_ (.A(_04283_),
    .B(_02365_),
    .Y(_04284_));
 sky130_fd_sc_hd__a211o_1 _10379_ (.A1(_04283_),
    .A2(\Oset[3][9] ),
    .B1(_03761_),
    .C1(_04284_),
    .X(_04285_));
 sky130_fd_sc_hd__nor2_1 _10380_ (.A(_04283_),
    .B(_02368_),
    .Y(_04286_));
 sky130_fd_sc_hd__a211o_1 _10381_ (.A1(_04283_),
    .A2(\Oset[1][9] ),
    .B1(_03764_),
    .C1(_04286_),
    .X(_04287_));
 sky130_fd_sc_hd__nand2_2 _10382_ (.A(_04285_),
    .B(_04287_),
    .Y(_04288_));
 sky130_fd_sc_hd__nand2_1 _10383_ (.A(_02363_),
    .B(_02163_),
    .Y(_04289_));
 sky130_fd_sc_hd__nor2_1 _10384_ (.A(_03760_),
    .B(_02357_),
    .Y(_04290_));
 sky130_fd_sc_hd__a211o_1 _10385_ (.A1(_03760_),
    .A2(\Qset[3][9] ),
    .B1(_03761_),
    .C1(_04290_),
    .X(_04291_));
 sky130_fd_sc_hd__nor2_1 _10386_ (.A(_03760_),
    .B(_02360_),
    .Y(_04292_));
 sky130_fd_sc_hd__a211o_1 _10387_ (.A1(_03760_),
    .A2(\Qset[1][9] ),
    .B1(_03764_),
    .C1(_04292_),
    .X(_04293_));
 sky130_fd_sc_hd__nand2_2 _10388_ (.A(_04291_),
    .B(_04293_),
    .Y(_04294_));
 sky130_fd_sc_hd__nand2_1 _10389_ (.A(_04294_),
    .B(_00582_),
    .Y(_04295_));
 sky130_fd_sc_hd__nand3_1 _10390_ (.A(_04289_),
    .B(_04295_),
    .C(_03770_),
    .Y(_04296_));
 sky130_fd_sc_hd__o21ai_1 _10391_ (.A1(_03770_),
    .A2(_04288_),
    .B1(_04296_),
    .Y(_04297_));
 sky130_fd_sc_hd__nand2_1 _10392_ (.A(_04297_),
    .B(_01156_),
    .Y(_04298_));
 sky130_fd_sc_hd__or2_1 _10393_ (.A(_01156_),
    .B(_02371_),
    .X(_04299_));
 sky130_fd_sc_hd__mux2_1 _10394_ (.A0(\H[2][9] ),
    .A1(\H[3][9] ),
    .S(_04282_),
    .X(_04300_));
 sky130_fd_sc_hd__nor2_1 _10395_ (.A(_04283_),
    .B(\H[0][9] ),
    .Y(_04301_));
 sky130_fd_sc_hd__buf_4 _10396_ (.A(_03773_),
    .X(_04302_));
 sky130_fd_sc_hd__clkbuf_4 _10397_ (.A(_03761_),
    .X(_04303_));
 sky130_fd_sc_hd__o21ai_1 _10398_ (.A1(\H[1][9] ),
    .A2(_04302_),
    .B1(_04303_),
    .Y(_04304_));
 sky130_fd_sc_hd__o2bb2a_1 _10399_ (.A1_N(_03764_),
    .A2_N(_04300_),
    .B1(_04301_),
    .B2(_04304_),
    .X(_04305_));
 sky130_fd_sc_hd__a21o_1 _10400_ (.A1(_04305_),
    .A2(_03768_),
    .B1(_00589_),
    .X(_04306_));
 sky130_fd_sc_hd__a31o_2 _10401_ (.A1(_04298_),
    .A2(_04299_),
    .A3(_03758_),
    .B1(_04306_),
    .X(_04307_));
 sky130_fd_sc_hd__nand2_8 _10402_ (.A(_04307_),
    .B(_02381_),
    .Y(_04308_));
 sky130_fd_sc_hd__clkinv_4 _10403_ (.A(_04308_),
    .Y(_04309_));
 sky130_fd_sc_hd__nor2_1 _10404_ (.A(_04281_),
    .B(_04309_),
    .Y(_04310_));
 sky130_fd_sc_hd__nand2_1 _10405_ (.A(_04280_),
    .B(_04310_),
    .Y(_04311_));
 sky130_fd_sc_hd__nand3b_1 _10406_ (.A_N(_04310_),
    .B(_04277_),
    .C(_04279_),
    .Y(_04312_));
 sky130_fd_sc_hd__nand3b_1 _10407_ (.A_N(_04263_),
    .B(_04311_),
    .C(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__nand2_1 _10408_ (.A(_04311_),
    .B(_04312_),
    .Y(_04314_));
 sky130_fd_sc_hd__nand2_1 _10409_ (.A(_04314_),
    .B(_04263_),
    .Y(_04315_));
 sky130_fd_sc_hd__nand2_1 _10410_ (.A(_04313_),
    .B(_04315_),
    .Y(_04316_));
 sky130_fd_sc_hd__inv_2 _10411_ (.A(_04316_),
    .Y(_04317_));
 sky130_fd_sc_hd__nand2_2 _10412_ (.A(_04262_),
    .B(_04317_),
    .Y(_04318_));
 sky130_fd_sc_hd__nand3_1 _10413_ (.A(_04234_),
    .B(_04261_),
    .C(_04316_),
    .Y(_04319_));
 sky130_fd_sc_hd__nand2_1 _10414_ (.A(_04318_),
    .B(_04319_),
    .Y(_04320_));
 sky130_fd_sc_hd__inv_2 _10415_ (.A(_03411_),
    .Y(_04321_));
 sky130_fd_sc_hd__nand2_1 _10416_ (.A(_04320_),
    .B(_04321_),
    .Y(_04322_));
 sky130_fd_sc_hd__nand3_1 _10417_ (.A(_04318_),
    .B(_03411_),
    .C(_04319_),
    .Y(_04323_));
 sky130_fd_sc_hd__nand2_1 _10418_ (.A(_04322_),
    .B(_04323_),
    .Y(_04324_));
 sky130_fd_sc_hd__nand2_1 _10419_ (.A(_04260_),
    .B(_04324_),
    .Y(_04325_));
 sky130_fd_sc_hd__inv_2 _10420_ (.A(_04324_),
    .Y(_04326_));
 sky130_fd_sc_hd__nand3_1 _10421_ (.A(_04244_),
    .B(_04326_),
    .C(_04239_),
    .Y(_04327_));
 sky130_fd_sc_hd__nand2_1 _10422_ (.A(_04325_),
    .B(_04327_),
    .Y(_04328_));
 sky130_fd_sc_hd__a32o_1 _10423_ (.A1(_03859_),
    .A2(_02620_),
    .A3(_03745_),
    .B1(_03835_),
    .B2(_03908_),
    .X(_04329_));
 sky130_fd_sc_hd__inv_2 _10424_ (.A(_04329_),
    .Y(_04330_));
 sky130_fd_sc_hd__nor2_1 _10425_ (.A(_03950_),
    .B(_04330_),
    .Y(_04331_));
 sky130_fd_sc_hd__inv_2 _10426_ (.A(_04331_),
    .Y(_04332_));
 sky130_fd_sc_hd__nand2_1 _10427_ (.A(_04328_),
    .B(_04332_),
    .Y(_04333_));
 sky130_fd_sc_hd__nand3_1 _10428_ (.A(_04325_),
    .B(_04327_),
    .C(_04331_),
    .Y(_04334_));
 sky130_fd_sc_hd__a21o_1 _10429_ (.A1(_04333_),
    .A2(_04334_),
    .B1(_04246_),
    .X(_04335_));
 sky130_fd_sc_hd__nand3_1 _10430_ (.A(_04333_),
    .B(_04246_),
    .C(_04334_),
    .Y(_04336_));
 sky130_fd_sc_hd__nand2_1 _10431_ (.A(_04335_),
    .B(_04336_),
    .Y(_04337_));
 sky130_fd_sc_hd__nand2_1 _10432_ (.A(_04337_),
    .B(_03746_),
    .Y(_04338_));
 sky130_fd_sc_hd__nand2_1 _10433_ (.A(_04194_),
    .B(_04157_),
    .Y(_04339_));
 sky130_fd_sc_hd__nand2_1 _10434_ (.A(_04040_),
    .B(_04028_),
    .Y(_04340_));
 sky130_fd_sc_hd__and2_1 _10435_ (.A(_04024_),
    .B(_04021_),
    .X(_04341_));
 sky130_fd_sc_hd__nor2_1 _10436_ (.A(_03899_),
    .B(_04309_),
    .Y(_04342_));
 sky130_fd_sc_hd__inv_2 _10437_ (.A(_04342_),
    .Y(_04343_));
 sky130_fd_sc_hd__and2_1 _10438_ (.A(_04018_),
    .B(_04014_),
    .X(_04344_));
 sky130_fd_sc_hd__inv_2 _10439_ (.A(_03859_),
    .Y(_04345_));
 sky130_fd_sc_hd__nor2_1 _10440_ (.A(_04345_),
    .B(_04025_),
    .Y(_04346_));
 sky130_fd_sc_hd__nand2_1 _10441_ (.A(_03652_),
    .B(_03868_),
    .Y(_04347_));
 sky130_fd_sc_hd__nand2_1 _10442_ (.A(_03652_),
    .B(_03876_),
    .Y(_04348_));
 sky130_fd_sc_hd__nand2_1 _10443_ (.A(_03506_),
    .B(_03868_),
    .Y(_04349_));
 sky130_fd_sc_hd__nand2_1 _10444_ (.A(_04348_),
    .B(_04349_),
    .Y(_04350_));
 sky130_fd_sc_hd__o21a_1 _10445_ (.A1(_04013_),
    .A2(_04347_),
    .B1(_04350_),
    .X(_04351_));
 sky130_fd_sc_hd__or2_1 _10446_ (.A(_04346_),
    .B(_04351_),
    .X(_04352_));
 sky130_fd_sc_hd__nand2_1 _10447_ (.A(_04351_),
    .B(_04346_),
    .Y(_04353_));
 sky130_fd_sc_hd__nand2_1 _10448_ (.A(_04352_),
    .B(_04353_),
    .Y(_04354_));
 sky130_fd_sc_hd__or2_1 _10449_ (.A(_04344_),
    .B(_04354_),
    .X(_04355_));
 sky130_fd_sc_hd__nand2_1 _10450_ (.A(_04354_),
    .B(_04344_),
    .Y(_04356_));
 sky130_fd_sc_hd__nand2_1 _10451_ (.A(_04355_),
    .B(_04356_),
    .Y(_04357_));
 sky130_fd_sc_hd__or2_1 _10452_ (.A(_04343_),
    .B(_04357_),
    .X(_04358_));
 sky130_fd_sc_hd__nand2_1 _10453_ (.A(_04357_),
    .B(_04343_),
    .Y(_04359_));
 sky130_fd_sc_hd__nand3b_1 _10454_ (.A_N(_04341_),
    .B(_04358_),
    .C(_04359_),
    .Y(_04360_));
 sky130_fd_sc_hd__nand2_1 _10455_ (.A(_04358_),
    .B(_04359_),
    .Y(_04361_));
 sky130_fd_sc_hd__nand2_1 _10456_ (.A(_04361_),
    .B(_04341_),
    .Y(_04362_));
 sky130_fd_sc_hd__nand2_1 _10457_ (.A(_04360_),
    .B(_04362_),
    .Y(_04363_));
 sky130_fd_sc_hd__nand2_1 _10458_ (.A(_04340_),
    .B(_04363_),
    .Y(_04364_));
 sky130_fd_sc_hd__inv_2 _10459_ (.A(_04363_),
    .Y(_04365_));
 sky130_fd_sc_hd__nand3_1 _10460_ (.A(_04040_),
    .B(_04365_),
    .C(_04028_),
    .Y(_04366_));
 sky130_fd_sc_hd__o21bai_1 _10461_ (.A1(_04151_),
    .A2(_04140_),
    .B1_N(_04138_),
    .Y(_04367_));
 sky130_fd_sc_hd__nor2_1 _10462_ (.A(_03205_),
    .B(_04050_),
    .Y(_04368_));
 sky130_fd_sc_hd__nand2_1 _10463_ (.A(_04074_),
    .B(_02963_),
    .Y(_04369_));
 sky130_fd_sc_hd__xor2_1 _10464_ (.A(_04369_),
    .B(_04124_),
    .X(_04370_));
 sky130_fd_sc_hd__or2_1 _10465_ (.A(_04368_),
    .B(_04370_),
    .X(_04371_));
 sky130_fd_sc_hd__nand2_1 _10466_ (.A(_04370_),
    .B(_04368_),
    .Y(_04372_));
 sky130_fd_sc_hd__nand2_1 _10467_ (.A(_04371_),
    .B(_04372_),
    .Y(_04373_));
 sky130_fd_sc_hd__nor2_1 _10468_ (.A(_04125_),
    .B(_04097_),
    .Y(_04374_));
 sky130_fd_sc_hd__inv_2 _10469_ (.A(_04129_),
    .Y(_04375_));
 sky130_fd_sc_hd__nor2_1 _10470_ (.A(_04374_),
    .B(_04375_),
    .Y(_04376_));
 sky130_fd_sc_hd__inv_2 _10471_ (.A(_04376_),
    .Y(_04377_));
 sky130_fd_sc_hd__or2_1 _10472_ (.A(_04373_),
    .B(_04377_),
    .X(_04378_));
 sky130_fd_sc_hd__nand2_1 _10473_ (.A(_04377_),
    .B(_04373_),
    .Y(_04379_));
 sky130_fd_sc_hd__nor2_1 _10474_ (.A(_03350_),
    .B(_04110_),
    .Y(_04380_));
 sky130_fd_sc_hd__a21bo_1 _10475_ (.A1(_04378_),
    .A2(_04379_),
    .B1_N(_04380_),
    .X(_04381_));
 sky130_fd_sc_hd__nand3b_1 _10476_ (.A_N(_04380_),
    .B(_04378_),
    .C(_04379_),
    .Y(_04382_));
 sky130_fd_sc_hd__nand2_1 _10477_ (.A(_04381_),
    .B(_04382_),
    .Y(_04383_));
 sky130_fd_sc_hd__a21oi_1 _10478_ (.A1(_04132_),
    .A2(_04134_),
    .B1(_04131_),
    .Y(_04384_));
 sky130_fd_sc_hd__nand2_1 _10479_ (.A(_04383_),
    .B(_04384_),
    .Y(_04385_));
 sky130_fd_sc_hd__or2_1 _10480_ (.A(_04384_),
    .B(_04383_),
    .X(_04386_));
 sky130_fd_sc_hd__nand3_1 _10481_ (.A(_04367_),
    .B(_04385_),
    .C(_04386_),
    .Y(_04387_));
 sky130_fd_sc_hd__nand2_1 _10482_ (.A(_04386_),
    .B(_04385_),
    .Y(_04388_));
 sky130_fd_sc_hd__a21oi_1 _10483_ (.A1(_04153_),
    .A2(_04139_),
    .B1(_04138_),
    .Y(_04389_));
 sky130_fd_sc_hd__nand2_1 _10484_ (.A(_04388_),
    .B(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hd__nand2_1 _10485_ (.A(_04387_),
    .B(_04390_),
    .Y(_04391_));
 sky130_fd_sc_hd__nand3_1 _10486_ (.A(_04364_),
    .B(_04366_),
    .C(_04391_),
    .Y(_04392_));
 sky130_fd_sc_hd__nand2_1 _10487_ (.A(_04340_),
    .B(_04365_),
    .Y(_04393_));
 sky130_fd_sc_hd__nand3_1 _10488_ (.A(_04040_),
    .B(_04028_),
    .C(_04363_),
    .Y(_04394_));
 sky130_fd_sc_hd__inv_2 _10489_ (.A(_04391_),
    .Y(_04395_));
 sky130_fd_sc_hd__nand3_1 _10490_ (.A(_04393_),
    .B(_04394_),
    .C(_04395_),
    .Y(_04396_));
 sky130_fd_sc_hd__nand2_1 _10491_ (.A(_04392_),
    .B(_04396_),
    .Y(_04397_));
 sky130_fd_sc_hd__inv_2 _10492_ (.A(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__nand2_1 _10493_ (.A(_04339_),
    .B(_04398_),
    .Y(_04399_));
 sky130_fd_sc_hd__nand3_1 _10494_ (.A(_04194_),
    .B(_04157_),
    .C(_04397_),
    .Y(_04400_));
 sky130_fd_sc_hd__nand3_1 _10495_ (.A(_04399_),
    .B(_03048_),
    .C(_04400_),
    .Y(_04401_));
 sky130_fd_sc_hd__a21o_1 _10496_ (.A1(_04364_),
    .A2(_04366_),
    .B1(_03048_),
    .X(_04402_));
 sky130_fd_sc_hd__nand3_1 _10497_ (.A(_04401_),
    .B(_04196_),
    .C(_04402_),
    .Y(_04403_));
 sky130_fd_sc_hd__nand3_1 _10498_ (.A(_04338_),
    .B(_00710_),
    .C(_04403_),
    .Y(_04404_));
 sky130_fd_sc_hd__nand2_1 _10499_ (.A(_03859_),
    .B(_02096_),
    .Y(_04405_));
 sky130_fd_sc_hd__nand3_1 _10500_ (.A(_04404_),
    .B(_00831_),
    .C(_04405_),
    .Y(_04406_));
 sky130_fd_sc_hd__nand2_1 _10501_ (.A(_04401_),
    .B(_04402_),
    .Y(_04407_));
 sky130_fd_sc_hd__nand2_1 _10502_ (.A(_04407_),
    .B(_04196_),
    .Y(_04408_));
 sky130_fd_sc_hd__nand3_1 _10503_ (.A(_04335_),
    .B(_03746_),
    .C(_04336_),
    .Y(_04409_));
 sky130_fd_sc_hd__nand3_1 _10504_ (.A(_04408_),
    .B(_04409_),
    .C(_00710_),
    .Y(_04410_));
 sky130_fd_sc_hd__nand2_1 _10505_ (.A(_04345_),
    .B(_02096_),
    .Y(_04411_));
 sky130_fd_sc_hd__nand3_1 _10506_ (.A(_04410_),
    .B(_02092_),
    .C(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__nand2_1 _10507_ (.A(_04406_),
    .B(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__clkbuf_4 _10508_ (.A(_03023_),
    .X(_04414_));
 sky130_fd_sc_hd__clkbuf_4 _10509_ (.A(_04414_),
    .X(_04415_));
 sky130_fd_sc_hd__a21o_1 _10510_ (.A1(\H[3][9] ),
    .A2(_03792_),
    .B1(_03794_),
    .X(_04416_));
 sky130_fd_sc_hd__a21o_1 _10511_ (.A1(\H[2][9] ),
    .A2(_04415_),
    .B1(_04416_),
    .X(_04417_));
 sky130_fd_sc_hd__a21oi_1 _10512_ (.A1(_04415_),
    .A2(\H[0][9] ),
    .B1(_03798_),
    .Y(_04418_));
 sky130_fd_sc_hd__o21ai_1 _10513_ (.A1(_02377_),
    .A2(_04415_),
    .B1(_04418_),
    .Y(_04419_));
 sky130_fd_sc_hd__a21oi_1 _10514_ (.A1(\Qset[3][9] ),
    .A2(_03791_),
    .B1(_03794_),
    .Y(_04420_));
 sky130_fd_sc_hd__nand2_1 _10515_ (.A(_04414_),
    .B(\Qset[2][9] ),
    .Y(_04421_));
 sky130_fd_sc_hd__a21oi_1 _10516_ (.A1(_04414_),
    .A2(\Qset[0][9] ),
    .B1(_03798_),
    .Y(_04422_));
 sky130_fd_sc_hd__nand2_1 _10517_ (.A(\Qset[1][9] ),
    .B(_03792_),
    .Y(_04423_));
 sky130_fd_sc_hd__a221o_1 _10518_ (.A1(_04420_),
    .A2(_04421_),
    .B1(_04422_),
    .B2(_04423_),
    .C1(_00621_),
    .X(_04424_));
 sky130_fd_sc_hd__a21oi_1 _10519_ (.A1(\Oset[3][9] ),
    .A2(_03791_),
    .B1(_03794_),
    .Y(_04425_));
 sky130_fd_sc_hd__nand2_1 _10520_ (.A(_04414_),
    .B(\Oset[2][9] ),
    .Y(_04426_));
 sky130_fd_sc_hd__a21oi_1 _10521_ (.A1(_04414_),
    .A2(\Oset[0][9] ),
    .B1(_03798_),
    .Y(_04427_));
 sky130_fd_sc_hd__nand2_1 _10522_ (.A(\Oset[1][9] ),
    .B(_03792_),
    .Y(_04428_));
 sky130_fd_sc_hd__a221o_1 _10523_ (.A1(_04425_),
    .A2(_04426_),
    .B1(_04427_),
    .B2(_04428_),
    .C1(_00647_),
    .X(_04429_));
 sky130_fd_sc_hd__a21oi_1 _10524_ (.A1(_04424_),
    .A2(_04429_),
    .B1(_01537_),
    .Y(_04430_));
 sky130_fd_sc_hd__a311o_2 _10525_ (.A1(_01537_),
    .A2(_04417_),
    .A3(_04419_),
    .B1(_00556_),
    .C1(_04430_),
    .X(_04431_));
 sky130_fd_sc_hd__o21ai_1 _10526_ (.A1(_00710_),
    .A2(_04308_),
    .B1(_04431_),
    .Y(_04432_));
 sky130_fd_sc_hd__nand2_1 _10527_ (.A(_04413_),
    .B(_04432_),
    .Y(_04433_));
 sky130_fd_sc_hd__nand3b_1 _10528_ (.A_N(_04432_),
    .B(_04406_),
    .C(_04412_),
    .Y(_04434_));
 sky130_fd_sc_hd__nand2_1 _10529_ (.A(_04433_),
    .B(_04434_),
    .Y(_04435_));
 sky130_fd_sc_hd__nor2_1 _10530_ (.A(_03752_),
    .B(_03755_),
    .Y(_04436_));
 sky130_fd_sc_hd__a21oi_1 _10531_ (.A1(_03756_),
    .A2(_03813_),
    .B1(_04436_),
    .Y(_04437_));
 sky130_fd_sc_hd__nor2_1 _10532_ (.A(_04435_),
    .B(_04437_),
    .Y(_04438_));
 sky130_fd_sc_hd__nand2_1 _10533_ (.A(_04437_),
    .B(_04435_),
    .Y(_04439_));
 sky130_fd_sc_hd__inv_2 _10534_ (.A(_04439_),
    .Y(_04440_));
 sky130_fd_sc_hd__nor2_1 _10535_ (.A(_04438_),
    .B(_04440_),
    .Y(_04441_));
 sky130_fd_sc_hd__or2_1 _10536_ (.A(_04255_),
    .B(_04441_),
    .X(_04442_));
 sky130_fd_sc_hd__nand2_1 _10537_ (.A(_04441_),
    .B(_04255_),
    .Y(_04443_));
 sky130_fd_sc_hd__nand2_2 _10538_ (.A(_04442_),
    .B(_04443_),
    .Y(_04444_));
 sky130_fd_sc_hd__nor2_1 _10539_ (.A(_02653_),
    .B(_04444_),
    .Y(_04445_));
 sky130_fd_sc_hd__a211o_1 _10540_ (.A1(_00933_),
    .A2(_02654_),
    .B1(_02753_),
    .C1(_04445_),
    .X(_04446_));
 sky130_fd_sc_hd__inv_2 _10541_ (.A(_04446_),
    .Y(_00253_));
 sky130_fd_sc_hd__nand2_1 _10542_ (.A(_04336_),
    .B(_04334_),
    .Y(_04447_));
 sky130_fd_sc_hd__inv_2 _10543_ (.A(_04447_),
    .Y(_04448_));
 sky130_fd_sc_hd__nand3_1 _10544_ (.A(_04241_),
    .B(_04240_),
    .C(_04324_),
    .Y(_04449_));
 sky130_fd_sc_hd__nand2_1 _10545_ (.A(_04320_),
    .B(_03411_),
    .Y(_04450_));
 sky130_fd_sc_hd__inv_2 _10546_ (.A(_04239_),
    .Y(_04451_));
 sky130_fd_sc_hd__nand3_1 _10547_ (.A(_04318_),
    .B(_04321_),
    .C(_04319_),
    .Y(_04452_));
 sky130_fd_sc_hd__a21boi_1 _10548_ (.A1(_04450_),
    .A2(_04451_),
    .B1_N(_04452_),
    .Y(_04453_));
 sky130_fd_sc_hd__nand2_1 _10549_ (.A(_04449_),
    .B(_04453_),
    .Y(_04454_));
 sky130_fd_sc_hd__nand2_1 _10550_ (.A(_04318_),
    .B(_04313_),
    .Y(_04455_));
 sky130_fd_sc_hd__or2_1 _10551_ (.A(_04278_),
    .B(_04276_),
    .X(_04456_));
 sky130_fd_sc_hd__and2_1 _10552_ (.A(_04311_),
    .B(_04456_),
    .X(_04457_));
 sky130_fd_sc_hd__inv_2 _10553_ (.A(_04270_),
    .Y(_04458_));
 sky130_fd_sc_hd__nor2_1 _10554_ (.A(_04458_),
    .B(_04309_),
    .Y(_04459_));
 sky130_fd_sc_hd__nor2_1 _10555_ (.A(_03897_),
    .B(_02897_),
    .Y(_04460_));
 sky130_fd_sc_hd__nand2_1 _10556_ (.A(_03790_),
    .B(_04460_),
    .Y(_04461_));
 sky130_fd_sc_hd__xor2_1 _10557_ (.A(_04265_),
    .B(_04461_),
    .X(_04462_));
 sky130_fd_sc_hd__or2_1 _10558_ (.A(_04459_),
    .B(_04462_),
    .X(_04463_));
 sky130_fd_sc_hd__nand2_1 _10559_ (.A(_04462_),
    .B(_04459_),
    .Y(_04464_));
 sky130_fd_sc_hd__nand2_1 _10560_ (.A(_04463_),
    .B(_04464_),
    .Y(_04465_));
 sky130_fd_sc_hd__inv_2 _10561_ (.A(_04275_),
    .Y(_04466_));
 sky130_fd_sc_hd__nor2_1 _10562_ (.A(_04266_),
    .B(_04466_),
    .Y(_04467_));
 sky130_fd_sc_hd__nand2_1 _10563_ (.A(_04465_),
    .B(_04467_),
    .Y(_04468_));
 sky130_fd_sc_hd__inv_2 _10564_ (.A(_04467_),
    .Y(_04469_));
 sky130_fd_sc_hd__nand3_1 _10565_ (.A(_04463_),
    .B(_04469_),
    .C(_04464_),
    .Y(_04470_));
 sky130_fd_sc_hd__nand2_1 _10566_ (.A(_02395_),
    .B(_02162_),
    .Y(_04471_));
 sky130_fd_sc_hd__inv_2 _10567_ (.A(\Qset[2][10] ),
    .Y(_04472_));
 sky130_fd_sc_hd__nor2_1 _10568_ (.A(_03759_),
    .B(_04472_),
    .Y(_04473_));
 sky130_fd_sc_hd__a211o_1 _10569_ (.A1(_04282_),
    .A2(\Qset[3][10] ),
    .B1(_03761_),
    .C1(_04473_),
    .X(_04474_));
 sky130_fd_sc_hd__nor2_1 _10570_ (.A(_03759_),
    .B(_02391_),
    .Y(_04475_));
 sky130_fd_sc_hd__a211o_1 _10571_ (.A1(_04282_),
    .A2(\Qset[1][10] ),
    .B1(_03345_),
    .C1(_04475_),
    .X(_04476_));
 sky130_fd_sc_hd__nand2_1 _10572_ (.A(_04474_),
    .B(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hd__nand2_1 _10573_ (.A(_04477_),
    .B(_00582_),
    .Y(_04478_));
 sky130_fd_sc_hd__nor2_1 _10574_ (.A(\Oset[3][10] ),
    .B(_03773_),
    .Y(_04479_));
 sky130_fd_sc_hd__o21ai_1 _10575_ (.A1(_04282_),
    .A2(\Oset[2][10] ),
    .B1(_03345_),
    .Y(_04480_));
 sky130_fd_sc_hd__nor2_1 _10576_ (.A(_04282_),
    .B(\Oset[0][10] ),
    .Y(_04481_));
 sky130_fd_sc_hd__o21ai_1 _10577_ (.A1(\Oset[1][10] ),
    .A2(_03773_),
    .B1(_03761_),
    .Y(_04482_));
 sky130_fd_sc_hd__o22a_2 _10578_ (.A1(_04479_),
    .A2(_04480_),
    .B1(_04481_),
    .B2(_04482_),
    .X(_04483_));
 sky130_fd_sc_hd__o21ai_1 _10579_ (.A1(_03770_),
    .A2(_04483_),
    .B1(_01156_),
    .Y(_04484_));
 sky130_fd_sc_hd__a31o_1 _10580_ (.A1(_04471_),
    .A2(_03770_),
    .A3(_04478_),
    .B1(_04484_),
    .X(_04485_));
 sky130_fd_sc_hd__nand2_1 _10581_ (.A(_02390_),
    .B(_00585_),
    .Y(_04486_));
 sky130_fd_sc_hd__mux2_1 _10582_ (.A0(\H[2][10] ),
    .A1(\H[3][10] ),
    .S(_04282_),
    .X(_04487_));
 sky130_fd_sc_hd__nor2_1 _10583_ (.A(_04283_),
    .B(\H[0][10] ),
    .Y(_04488_));
 sky130_fd_sc_hd__o21ai_1 _10584_ (.A1(\H[1][10] ),
    .A2(_04302_),
    .B1(_03761_),
    .Y(_04489_));
 sky130_fd_sc_hd__o2bb2a_1 _10585_ (.A1_N(_03764_),
    .A2_N(_04487_),
    .B1(_04488_),
    .B2(_04489_),
    .X(_04490_));
 sky130_fd_sc_hd__nor2_1 _10586_ (.A(_03758_),
    .B(_04490_),
    .Y(_04491_));
 sky130_fd_sc_hd__a31o_1 _10587_ (.A1(_04485_),
    .A2(_03758_),
    .A3(_04486_),
    .B1(_04491_),
    .X(_04492_));
 sky130_fd_sc_hd__nand2_2 _10588_ (.A(_04492_),
    .B(_01553_),
    .Y(_04493_));
 sky130_fd_sc_hd__nand2_8 _10589_ (.A(_04493_),
    .B(_02403_),
    .Y(_04494_));
 sky130_fd_sc_hd__inv_2 _10590_ (.A(_04494_),
    .Y(_04495_));
 sky130_fd_sc_hd__nor2_1 _10591_ (.A(_04281_),
    .B(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__nand3_1 _10592_ (.A(_04468_),
    .B(_04470_),
    .C(_04496_),
    .Y(_04497_));
 sky130_fd_sc_hd__nand2_1 _10593_ (.A(_04465_),
    .B(_04469_),
    .Y(_04498_));
 sky130_fd_sc_hd__inv_2 _10594_ (.A(_04496_),
    .Y(_04499_));
 sky130_fd_sc_hd__nand3_1 _10595_ (.A(_04463_),
    .B(_04467_),
    .C(_04464_),
    .Y(_04500_));
 sky130_fd_sc_hd__nand3_1 _10596_ (.A(_04498_),
    .B(_04499_),
    .C(_04500_),
    .Y(_04501_));
 sky130_fd_sc_hd__nand3b_2 _10597_ (.A_N(_04457_),
    .B(_04497_),
    .C(_04501_),
    .Y(_04502_));
 sky130_fd_sc_hd__nand2_1 _10598_ (.A(_04497_),
    .B(_04501_),
    .Y(_04503_));
 sky130_fd_sc_hd__nand2_1 _10599_ (.A(_04503_),
    .B(_04457_),
    .Y(_04504_));
 sky130_fd_sc_hd__nand2_1 _10600_ (.A(_04502_),
    .B(_04504_),
    .Y(_04505_));
 sky130_fd_sc_hd__inv_2 _10601_ (.A(_04505_),
    .Y(_04506_));
 sky130_fd_sc_hd__nand2_1 _10602_ (.A(_04455_),
    .B(_04506_),
    .Y(_04507_));
 sky130_fd_sc_hd__nand3_1 _10603_ (.A(_04318_),
    .B(_04505_),
    .C(_04313_),
    .Y(_04508_));
 sky130_fd_sc_hd__nand2_1 _10604_ (.A(_04507_),
    .B(_04508_),
    .Y(_04509_));
 sky130_fd_sc_hd__nand2_1 _10605_ (.A(_04509_),
    .B(_03564_),
    .Y(_04510_));
 sky130_fd_sc_hd__nand3b_1 _10606_ (.A_N(_03564_),
    .B(_04507_),
    .C(_04508_),
    .Y(_04511_));
 sky130_fd_sc_hd__nand2_1 _10607_ (.A(_04510_),
    .B(_04511_),
    .Y(_04512_));
 sky130_fd_sc_hd__inv_2 _10608_ (.A(_04512_),
    .Y(_04513_));
 sky130_fd_sc_hd__nand2_1 _10609_ (.A(_04454_),
    .B(_04513_),
    .Y(_04514_));
 sky130_fd_sc_hd__nand3_1 _10610_ (.A(_04512_),
    .B(_04449_),
    .C(_04453_),
    .Y(_04515_));
 sky130_fd_sc_hd__nand2_1 _10611_ (.A(_04514_),
    .B(_04515_),
    .Y(_04516_));
 sky130_fd_sc_hd__inv_2 _10612_ (.A(_04516_),
    .Y(_04517_));
 sky130_fd_sc_hd__or2_1 _10613_ (.A(_03950_),
    .B(_03948_),
    .X(_04518_));
 sky130_fd_sc_hd__nand2_1 _10614_ (.A(_04518_),
    .B(_03951_),
    .Y(_04519_));
 sky130_fd_sc_hd__nand2_1 _10615_ (.A(_04517_),
    .B(_04519_),
    .Y(_04520_));
 sky130_fd_sc_hd__inv_2 _10616_ (.A(_04519_),
    .Y(_04521_));
 sky130_fd_sc_hd__nand2_1 _10617_ (.A(_04516_),
    .B(_04521_),
    .Y(_04522_));
 sky130_fd_sc_hd__nand2_1 _10618_ (.A(_04520_),
    .B(_04522_),
    .Y(_04523_));
 sky130_fd_sc_hd__inv_2 _10619_ (.A(_04523_),
    .Y(_04524_));
 sky130_fd_sc_hd__nand2_1 _10620_ (.A(_04448_),
    .B(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__nand2_1 _10621_ (.A(_04447_),
    .B(_04523_),
    .Y(_04526_));
 sky130_fd_sc_hd__nand3_2 _10622_ (.A(_04525_),
    .B(_03746_),
    .C(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__nand3_1 _10623_ (.A(_04398_),
    .B(_04192_),
    .C(_04159_),
    .Y(_04528_));
 sky130_fd_sc_hd__inv_2 _10624_ (.A(_04157_),
    .Y(_04529_));
 sky130_fd_sc_hd__a21boi_1 _10625_ (.A1(_04529_),
    .A2(_04392_),
    .B1_N(_04396_),
    .Y(_04530_));
 sky130_fd_sc_hd__nand2_1 _10626_ (.A(_04528_),
    .B(_04530_),
    .Y(_04531_));
 sky130_fd_sc_hd__nand2b_1 _10627_ (.A_N(_04040_),
    .B(_04365_),
    .Y(_04532_));
 sky130_fd_sc_hd__nor2_1 _10628_ (.A(_04011_),
    .B(_04027_),
    .Y(_04533_));
 sky130_fd_sc_hd__a21boi_1 _10629_ (.A1(_04533_),
    .A2(_04362_),
    .B1_N(_04360_),
    .Y(_04534_));
 sky130_fd_sc_hd__nand2_1 _10630_ (.A(_04532_),
    .B(_04534_),
    .Y(_04535_));
 sky130_fd_sc_hd__nor2_1 _10631_ (.A(_03899_),
    .B(_04495_),
    .Y(_04536_));
 sky130_fd_sc_hd__inv_2 _10632_ (.A(_04536_),
    .Y(_04537_));
 sky130_fd_sc_hd__o21a_1 _10633_ (.A1(_04349_),
    .A2(_04348_),
    .B1(_04353_),
    .X(_04538_));
 sky130_fd_sc_hd__nor2_1 _10634_ (.A(_04345_),
    .B(_04309_),
    .Y(_04539_));
 sky130_fd_sc_hd__inv_2 _10635_ (.A(_03874_),
    .Y(_04540_));
 sky130_fd_sc_hd__nor2_1 _10636_ (.A(_04105_),
    .B(_02387_),
    .Y(_04541_));
 sky130_fd_sc_hd__nand2_1 _10637_ (.A(_02567_),
    .B(\Oset[1][10] ),
    .Y(_04542_));
 sky130_fd_sc_hd__inv_2 _10638_ (.A(_04542_),
    .Y(_04543_));
 sky130_fd_sc_hd__nor2_1 _10639_ (.A(_02567_),
    .B(_02384_),
    .Y(_04544_));
 sky130_fd_sc_hd__a211o_1 _10640_ (.A1(_04105_),
    .A2(\Oset[3][10] ),
    .B1(_04045_),
    .C1(_04544_),
    .X(_04545_));
 sky130_fd_sc_hd__o31ai_4 _10641_ (.A1(_04042_),
    .A2(_04541_),
    .A3(_04543_),
    .B1(_04545_),
    .Y(_04546_));
 sky130_fd_sc_hd__a21oi_1 _10642_ (.A1(_04546_),
    .A2(_03781_),
    .B1(_00585_),
    .Y(_04547_));
 sky130_fd_sc_hd__nor2_1 _10643_ (.A(_04105_),
    .B(_04472_),
    .Y(_04548_));
 sky130_fd_sc_hd__a211o_1 _10644_ (.A1(_04105_),
    .A2(\Qset[3][10] ),
    .B1(_04045_),
    .C1(_04548_),
    .X(_04549_));
 sky130_fd_sc_hd__nor2_1 _10645_ (.A(_04105_),
    .B(_02391_),
    .Y(_04550_));
 sky130_fd_sc_hd__a211o_1 _10646_ (.A1(_04105_),
    .A2(\Qset[1][10] ),
    .B1(_04042_),
    .C1(_04550_),
    .X(_04551_));
 sky130_fd_sc_hd__nand2_2 _10647_ (.A(_04549_),
    .B(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__o21ai_1 _10648_ (.A1(_02163_),
    .A2(_04552_),
    .B1(_02796_),
    .Y(_04553_));
 sky130_fd_sc_hd__nand2_1 _10649_ (.A(_04547_),
    .B(_04553_),
    .Y(_04554_));
 sky130_fd_sc_hd__a221oi_4 _10650_ (.A1(_03768_),
    .A2(_04540_),
    .B1(_04554_),
    .B2(_02811_),
    .C1(_00589_),
    .Y(_04555_));
 sky130_fd_sc_hd__nand2_1 _10651_ (.A(_03790_),
    .B(_04555_),
    .Y(_04556_));
 sky130_fd_sc_hd__nor2_1 _10652_ (.A(_04347_),
    .B(_04556_),
    .Y(_04557_));
 sky130_fd_sc_hd__nand2_1 _10653_ (.A(_04556_),
    .B(_04347_),
    .Y(_04558_));
 sky130_fd_sc_hd__nor2b_1 _10654_ (.A(_04557_),
    .B_N(_04558_),
    .Y(_04559_));
 sky130_fd_sc_hd__xnor2_1 _10655_ (.A(_04539_),
    .B(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__or2_1 _10656_ (.A(_04538_),
    .B(_04560_),
    .X(_04561_));
 sky130_fd_sc_hd__nand2_1 _10657_ (.A(_04560_),
    .B(_04538_),
    .Y(_04562_));
 sky130_fd_sc_hd__nand2_1 _10658_ (.A(_04561_),
    .B(_04562_),
    .Y(_04563_));
 sky130_fd_sc_hd__or2_1 _10659_ (.A(_04537_),
    .B(_04563_),
    .X(_04564_));
 sky130_fd_sc_hd__nand2_1 _10660_ (.A(_04563_),
    .B(_04537_),
    .Y(_04565_));
 sky130_fd_sc_hd__nand2_1 _10661_ (.A(_04358_),
    .B(_04355_),
    .Y(_04566_));
 sky130_fd_sc_hd__a21o_1 _10662_ (.A1(_04564_),
    .A2(_04565_),
    .B1(_04566_),
    .X(_04567_));
 sky130_fd_sc_hd__nand3_2 _10663_ (.A(_04564_),
    .B(_04566_),
    .C(_04565_),
    .Y(_04568_));
 sky130_fd_sc_hd__nand2_1 _10664_ (.A(_04567_),
    .B(_04568_),
    .Y(_04569_));
 sky130_fd_sc_hd__inv_2 _10665_ (.A(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__nand2_2 _10666_ (.A(_04535_),
    .B(_04570_),
    .Y(_04571_));
 sky130_fd_sc_hd__nand3_1 _10667_ (.A(_04532_),
    .B(_04534_),
    .C(_04569_),
    .Y(_04572_));
 sky130_fd_sc_hd__nand2_1 _10668_ (.A(_04571_),
    .B(_04572_),
    .Y(_04573_));
 sky130_fd_sc_hd__nand2_1 _10669_ (.A(_04387_),
    .B(_04386_),
    .Y(_04574_));
 sky130_fd_sc_hd__nor2_1 _10670_ (.A(_03507_),
    .B(_04110_),
    .Y(_04575_));
 sky130_fd_sc_hd__o21a_1 _10671_ (.A1(_04124_),
    .A2(_04369_),
    .B1(_04372_),
    .X(_04576_));
 sky130_fd_sc_hd__nor2_1 _10672_ (.A(_03350_),
    .B(_04050_),
    .Y(_04577_));
 sky130_fd_sc_hd__nand2_1 _10673_ (.A(_04096_),
    .B(_03020_),
    .Y(_04578_));
 sky130_fd_sc_hd__nor2_1 _10674_ (.A(_04369_),
    .B(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hd__a22o_1 _10675_ (.A1(_04074_),
    .A2(_03020_),
    .B1(_04096_),
    .B2(_02963_),
    .X(_04580_));
 sky130_fd_sc_hd__and2b_1 _10676_ (.A_N(_04579_),
    .B(_04580_),
    .X(_04581_));
 sky130_fd_sc_hd__xnor2_1 _10677_ (.A(_04577_),
    .B(_04581_),
    .Y(_04582_));
 sky130_fd_sc_hd__nor2_1 _10678_ (.A(_04576_),
    .B(_04582_),
    .Y(_04583_));
 sky130_fd_sc_hd__nand2_1 _10679_ (.A(_04582_),
    .B(_04576_),
    .Y(_04584_));
 sky130_fd_sc_hd__and2b_1 _10680_ (.A_N(_04583_),
    .B(_04584_),
    .X(_04585_));
 sky130_fd_sc_hd__xnor2_1 _10681_ (.A(_04575_),
    .B(_04585_),
    .Y(_04586_));
 sky130_fd_sc_hd__o21a_1 _10682_ (.A1(_04376_),
    .A2(_04373_),
    .B1(_04381_),
    .X(_04587_));
 sky130_fd_sc_hd__nor2_1 _10683_ (.A(_04586_),
    .B(_04587_),
    .Y(_04588_));
 sky130_fd_sc_hd__inv_2 _10684_ (.A(_04588_),
    .Y(_04589_));
 sky130_fd_sc_hd__nand2_1 _10685_ (.A(_04587_),
    .B(_04586_),
    .Y(_04590_));
 sky130_fd_sc_hd__nand2_1 _10686_ (.A(_04589_),
    .B(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__inv_2 _10687_ (.A(_04591_),
    .Y(_04592_));
 sky130_fd_sc_hd__nand2_1 _10688_ (.A(_04574_),
    .B(_04592_),
    .Y(_04593_));
 sky130_fd_sc_hd__nand3_1 _10689_ (.A(_04591_),
    .B(_04387_),
    .C(_04386_),
    .Y(_04594_));
 sky130_fd_sc_hd__nand2_1 _10690_ (.A(_04593_),
    .B(_04594_),
    .Y(_04595_));
 sky130_fd_sc_hd__nand2_1 _10691_ (.A(_04573_),
    .B(_04595_),
    .Y(_04596_));
 sky130_fd_sc_hd__nand3b_1 _10692_ (.A_N(_04595_),
    .B(_04571_),
    .C(_04572_),
    .Y(_04597_));
 sky130_fd_sc_hd__nand2_1 _10693_ (.A(_04596_),
    .B(_04597_),
    .Y(_04598_));
 sky130_fd_sc_hd__inv_2 _10694_ (.A(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__nand2_1 _10695_ (.A(_04531_),
    .B(_04599_),
    .Y(_04600_));
 sky130_fd_sc_hd__nand3_1 _10696_ (.A(_04598_),
    .B(_04528_),
    .C(_04530_),
    .Y(_04601_));
 sky130_fd_sc_hd__nand2_1 _10697_ (.A(_04600_),
    .B(_04601_),
    .Y(_04602_));
 sky130_fd_sc_hd__nand2_1 _10698_ (.A(_04602_),
    .B(_03048_),
    .Y(_04603_));
 sky130_fd_sc_hd__a21oi_1 _10699_ (.A1(_04573_),
    .A2(_03751_),
    .B1(_03745_),
    .Y(_04604_));
 sky130_fd_sc_hd__nand2_1 _10700_ (.A(_04603_),
    .B(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__nand3_1 _10701_ (.A(_04527_),
    .B(_04605_),
    .C(_00710_),
    .Y(_04606_));
 sky130_fd_sc_hd__inv_2 _10702_ (.A(_04555_),
    .Y(_04607_));
 sky130_fd_sc_hd__nand2_1 _10703_ (.A(_04607_),
    .B(_02096_),
    .Y(_04608_));
 sky130_fd_sc_hd__nand2_1 _10704_ (.A(_04606_),
    .B(_04608_),
    .Y(_04609_));
 sky130_fd_sc_hd__nand2_1 _10705_ (.A(_04609_),
    .B(_00831_),
    .Y(_04610_));
 sky130_fd_sc_hd__nand3_1 _10706_ (.A(_04606_),
    .B(_02092_),
    .C(_04608_),
    .Y(_04611_));
 sky130_fd_sc_hd__nand2_1 _10707_ (.A(_04610_),
    .B(_04611_),
    .Y(_04612_));
 sky130_fd_sc_hd__a21o_1 _10708_ (.A1(\H[3][10] ),
    .A2(_03792_),
    .B1(_03794_),
    .X(_04613_));
 sky130_fd_sc_hd__a21o_1 _10709_ (.A1(\H[2][10] ),
    .A2(_04414_),
    .B1(_04613_),
    .X(_04614_));
 sky130_fd_sc_hd__a21oi_1 _10710_ (.A1(_04414_),
    .A2(\H[0][10] ),
    .B1(_03798_),
    .Y(_04615_));
 sky130_fd_sc_hd__o21ai_1 _10711_ (.A1(_02400_),
    .A2(_04415_),
    .B1(_04615_),
    .Y(_04616_));
 sky130_fd_sc_hd__nand2_1 _10712_ (.A(_03023_),
    .B(\Qset[0][10] ),
    .Y(_04617_));
 sky130_fd_sc_hd__nand2_1 _10713_ (.A(\Qset[1][10] ),
    .B(_03791_),
    .Y(_04618_));
 sky130_fd_sc_hd__a21oi_1 _10714_ (.A1(\Qset[3][10] ),
    .A2(_03791_),
    .B1(_03794_),
    .Y(_04619_));
 sky130_fd_sc_hd__nand2_1 _10715_ (.A(_03023_),
    .B(\Qset[2][10] ),
    .Y(_04620_));
 sky130_fd_sc_hd__a32o_1 _10716_ (.A1(_04617_),
    .A2(_04618_),
    .A3(_03794_),
    .B1(_04619_),
    .B2(_04620_),
    .X(_04621_));
 sky130_fd_sc_hd__nand2_1 _10717_ (.A(_03023_),
    .B(\Oset[0][10] ),
    .Y(_04622_));
 sky130_fd_sc_hd__nand2_1 _10718_ (.A(\Oset[1][10] ),
    .B(_03791_),
    .Y(_04623_));
 sky130_fd_sc_hd__a21oi_1 _10719_ (.A1(\Oset[3][10] ),
    .A2(_03791_),
    .B1(_03027_),
    .Y(_04624_));
 sky130_fd_sc_hd__nand2_1 _10720_ (.A(_03023_),
    .B(\Oset[2][10] ),
    .Y(_04625_));
 sky130_fd_sc_hd__a32o_1 _10721_ (.A1(_04622_),
    .A2(_04623_),
    .A3(_03794_),
    .B1(_04624_),
    .B2(_04625_),
    .X(_04626_));
 sky130_fd_sc_hd__mux2_1 _10722_ (.A0(_04621_),
    .A1(_04626_),
    .S(_00621_),
    .X(_04627_));
 sky130_fd_sc_hd__nor2_1 _10723_ (.A(_01537_),
    .B(_04627_),
    .Y(_04628_));
 sky130_fd_sc_hd__a311o_2 _10724_ (.A1(_01537_),
    .A2(_04614_),
    .A3(_04616_),
    .B1(_00556_),
    .C1(_04628_),
    .X(_04629_));
 sky130_fd_sc_hd__o21ai_2 _10725_ (.A1(_00624_),
    .A2(_04494_),
    .B1(_04629_),
    .Y(_04630_));
 sky130_fd_sc_hd__nand2_1 _10726_ (.A(_04612_),
    .B(_04630_),
    .Y(_04631_));
 sky130_fd_sc_hd__inv_2 _10727_ (.A(_04630_),
    .Y(_04632_));
 sky130_fd_sc_hd__nand3_2 _10728_ (.A(_04610_),
    .B(_04611_),
    .C(_04632_),
    .Y(_04633_));
 sky130_fd_sc_hd__nand2_1 _10729_ (.A(_04631_),
    .B(_04633_),
    .Y(_04634_));
 sky130_fd_sc_hd__nand2_1 _10730_ (.A(_04634_),
    .B(_04434_),
    .Y(_04635_));
 sky130_fd_sc_hd__nand3b_1 _10731_ (.A_N(_04434_),
    .B(_04631_),
    .C(_04633_),
    .Y(_04636_));
 sky130_fd_sc_hd__nand2_1 _10732_ (.A(_04635_),
    .B(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__inv_2 _10733_ (.A(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__o21bai_1 _10734_ (.A1(_04255_),
    .A2(_04440_),
    .B1_N(_04438_),
    .Y(_04639_));
 sky130_fd_sc_hd__or2_1 _10735_ (.A(_04638_),
    .B(_04639_),
    .X(_04640_));
 sky130_fd_sc_hd__nand2_1 _10736_ (.A(_04639_),
    .B(_04638_),
    .Y(_04641_));
 sky130_fd_sc_hd__and2_2 _10737_ (.A(_04640_),
    .B(_04641_),
    .X(_04642_));
 sky130_fd_sc_hd__nor2_1 _10738_ (.A(_02653_),
    .B(_04642_),
    .Y(_04643_));
 sky130_fd_sc_hd__a211o_1 _10739_ (.A1(_00959_),
    .A2(_02654_),
    .B1(_02753_),
    .C1(_04643_),
    .X(_04644_));
 sky130_fd_sc_hd__inv_2 _10740_ (.A(_04644_),
    .Y(_00254_));
 sky130_fd_sc_hd__nand2_1 _10741_ (.A(_04517_),
    .B(_04521_),
    .Y(_04645_));
 sky130_fd_sc_hd__nand2_1 _10742_ (.A(_04526_),
    .B(_04645_),
    .Y(_04646_));
 sky130_fd_sc_hd__nand2_1 _10743_ (.A(_04514_),
    .B(_04511_),
    .Y(_04647_));
 sky130_fd_sc_hd__nand2_1 _10744_ (.A(_03701_),
    .B(_03703_),
    .Y(_04648_));
 sky130_fd_sc_hd__nand2_1 _10745_ (.A(_04507_),
    .B(_04502_),
    .Y(_04649_));
 sky130_fd_sc_hd__nand2_1 _10746_ (.A(_04308_),
    .B(_04460_),
    .Y(_04650_));
 sky130_fd_sc_hd__nor2_1 _10747_ (.A(_03897_),
    .B(_02904_),
    .Y(_04651_));
 sky130_fd_sc_hd__nand2_1 _10748_ (.A(_03790_),
    .B(_04651_),
    .Y(_04652_));
 sky130_fd_sc_hd__nor2_1 _10749_ (.A(_04650_),
    .B(_04652_),
    .Y(_04653_));
 sky130_fd_sc_hd__nand2_1 _10750_ (.A(_04652_),
    .B(_04650_),
    .Y(_04654_));
 sky130_fd_sc_hd__inv_2 _10751_ (.A(_04654_),
    .Y(_04655_));
 sky130_fd_sc_hd__nand2_1 _10752_ (.A(_04494_),
    .B(_04270_),
    .Y(_04656_));
 sky130_fd_sc_hd__o21ai_1 _10753_ (.A1(_04653_),
    .A2(_04655_),
    .B1(_04656_),
    .Y(_04657_));
 sky130_fd_sc_hd__inv_2 _10754_ (.A(_04656_),
    .Y(_04658_));
 sky130_fd_sc_hd__nand3b_1 _10755_ (.A_N(_04653_),
    .B(_04658_),
    .C(_04654_),
    .Y(_04659_));
 sky130_fd_sc_hd__nand2_1 _10756_ (.A(_04657_),
    .B(_04659_),
    .Y(_04660_));
 sky130_fd_sc_hd__nand2_1 _10757_ (.A(_04461_),
    .B(_04265_),
    .Y(_04661_));
 sky130_fd_sc_hd__nor2_1 _10758_ (.A(_04265_),
    .B(_04461_),
    .Y(_04662_));
 sky130_fd_sc_hd__a21oi_2 _10759_ (.A1(_04661_),
    .A2(_04459_),
    .B1(_04662_),
    .Y(_04663_));
 sky130_fd_sc_hd__inv_2 _10760_ (.A(_04663_),
    .Y(_04664_));
 sky130_fd_sc_hd__nand2_1 _10761_ (.A(_04660_),
    .B(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hd__nand3_1 _10762_ (.A(_04657_),
    .B(_04659_),
    .C(_04663_),
    .Y(_04666_));
 sky130_fd_sc_hd__nand2_1 _10763_ (.A(_04665_),
    .B(_04666_),
    .Y(_04667_));
 sky130_fd_sc_hd__nand2_1 _10764_ (.A(_04302_),
    .B(_03861_),
    .Y(_04668_));
 sky130_fd_sc_hd__a21oi_1 _10765_ (.A1(_02423_),
    .A2(_04283_),
    .B1(_03764_),
    .Y(_04669_));
 sky130_fd_sc_hd__mux2_1 _10766_ (.A0(\H[2][11] ),
    .A1(\H[3][11] ),
    .S(_03760_),
    .X(_04670_));
 sky130_fd_sc_hd__a22o_1 _10767_ (.A1(_04668_),
    .A2(_04669_),
    .B1(_04670_),
    .B2(_03764_),
    .X(_04671_));
 sky130_fd_sc_hd__nand2_1 _10768_ (.A(_02412_),
    .B(_02162_),
    .Y(_04672_));
 sky130_fd_sc_hd__nor2_1 _10769_ (.A(_04282_),
    .B(_02406_),
    .Y(_04673_));
 sky130_fd_sc_hd__a211o_1 _10770_ (.A1(_04282_),
    .A2(\Qset[3][11] ),
    .B1(_03761_),
    .C1(_04673_),
    .X(_04674_));
 sky130_fd_sc_hd__nor2_1 _10771_ (.A(_03759_),
    .B(_02409_),
    .Y(_04675_));
 sky130_fd_sc_hd__a211o_1 _10772_ (.A1(_04282_),
    .A2(\Qset[1][11] ),
    .B1(_03345_),
    .C1(_04675_),
    .X(_04676_));
 sky130_fd_sc_hd__nand2_1 _10773_ (.A(_04674_),
    .B(_04676_),
    .Y(_04677_));
 sky130_fd_sc_hd__nand2_1 _10774_ (.A(_04677_),
    .B(_00582_),
    .Y(_04678_));
 sky130_fd_sc_hd__nor2_1 _10775_ (.A(\Oset[3][11] ),
    .B(_03341_),
    .Y(_04679_));
 sky130_fd_sc_hd__o21ai_1 _10776_ (.A1(_03498_),
    .A2(\Oset[2][11] ),
    .B1(_03345_),
    .Y(_04680_));
 sky130_fd_sc_hd__nor2_1 _10777_ (.A(_03759_),
    .B(\Oset[0][11] ),
    .Y(_04681_));
 sky130_fd_sc_hd__o21ai_1 _10778_ (.A1(\Oset[1][11] ),
    .A2(_03341_),
    .B1(_03004_),
    .Y(_04682_));
 sky130_fd_sc_hd__o22a_2 _10779_ (.A1(_04679_),
    .A2(_04680_),
    .B1(_04681_),
    .B2(_04682_),
    .X(_04683_));
 sky130_fd_sc_hd__nor2_1 _10780_ (.A(_02540_),
    .B(_04683_),
    .Y(_04684_));
 sky130_fd_sc_hd__or2_1 _10781_ (.A(_00584_),
    .B(_04684_),
    .X(_04685_));
 sky130_fd_sc_hd__a31o_1 _10782_ (.A1(_03770_),
    .A2(_04672_),
    .A3(_04678_),
    .B1(_04685_),
    .X(_04686_));
 sky130_fd_sc_hd__a21oi_1 _10783_ (.A1(_02419_),
    .A2(_00584_),
    .B1(_03768_),
    .Y(_04687_));
 sky130_fd_sc_hd__a22o_1 _10784_ (.A1(_03768_),
    .A2(_04671_),
    .B1(_04686_),
    .B2(_04687_),
    .X(_04688_));
 sky130_fd_sc_hd__nand2_2 _10785_ (.A(_04688_),
    .B(_01553_),
    .Y(_04689_));
 sky130_fd_sc_hd__nand2_8 _10786_ (.A(_04689_),
    .B(_02426_),
    .Y(_04690_));
 sky130_fd_sc_hd__inv_6 _10787_ (.A(_04690_),
    .Y(_04691_));
 sky130_fd_sc_hd__nor2_1 _10788_ (.A(_04281_),
    .B(_04691_),
    .Y(_04692_));
 sky130_fd_sc_hd__nand2_1 _10789_ (.A(_04667_),
    .B(_04692_),
    .Y(_04693_));
 sky130_fd_sc_hd__nand3b_1 _10790_ (.A_N(_04692_),
    .B(_04665_),
    .C(_04666_),
    .Y(_04694_));
 sky130_fd_sc_hd__nand2_2 _10791_ (.A(_04693_),
    .B(_04694_),
    .Y(_04695_));
 sky130_fd_sc_hd__a21boi_2 _10792_ (.A1(_04468_),
    .A2(_04496_),
    .B1_N(_04470_),
    .Y(_04696_));
 sky130_fd_sc_hd__xor2_2 _10793_ (.A(_04695_),
    .B(_04696_),
    .X(_04697_));
 sky130_fd_sc_hd__nand2_1 _10794_ (.A(_04649_),
    .B(_04697_),
    .Y(_04698_));
 sky130_fd_sc_hd__inv_2 _10795_ (.A(_04502_),
    .Y(_04699_));
 sky130_fd_sc_hd__nor2_1 _10796_ (.A(_04699_),
    .B(_04697_),
    .Y(_04700_));
 sky130_fd_sc_hd__nand2_1 _10797_ (.A(_04507_),
    .B(_04700_),
    .Y(_04701_));
 sky130_fd_sc_hd__nand3b_1 _10798_ (.A_N(_04648_),
    .B(_04698_),
    .C(_04701_),
    .Y(_04702_));
 sky130_fd_sc_hd__nand2_1 _10799_ (.A(_04697_),
    .B(_04699_),
    .Y(_04703_));
 sky130_fd_sc_hd__nand3_1 _10800_ (.A(_04455_),
    .B(_04506_),
    .C(_04697_),
    .Y(_04704_));
 sky130_fd_sc_hd__nand3_1 _10801_ (.A(_04701_),
    .B(_04703_),
    .C(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__nand2_1 _10802_ (.A(_04705_),
    .B(_04648_),
    .Y(_04706_));
 sky130_fd_sc_hd__nand2_1 _10803_ (.A(_04702_),
    .B(_04706_),
    .Y(_04707_));
 sky130_fd_sc_hd__inv_2 _10804_ (.A(_04707_),
    .Y(_04708_));
 sky130_fd_sc_hd__nand2_1 _10805_ (.A(_04647_),
    .B(_04708_),
    .Y(_04709_));
 sky130_fd_sc_hd__nand3_1 _10806_ (.A(_04514_),
    .B(_04707_),
    .C(_04511_),
    .Y(_04710_));
 sky130_fd_sc_hd__nand2_1 _10807_ (.A(_04709_),
    .B(_04710_),
    .Y(_04711_));
 sky130_fd_sc_hd__nand2_1 _10808_ (.A(_03955_),
    .B(_03951_),
    .Y(_04712_));
 sky130_fd_sc_hd__or2b_1 _10809_ (.A(_03956_),
    .B_N(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__nand2_1 _10810_ (.A(_04711_),
    .B(_04713_),
    .Y(_04714_));
 sky130_fd_sc_hd__inv_2 _10811_ (.A(_04713_),
    .Y(_04715_));
 sky130_fd_sc_hd__nand3_1 _10812_ (.A(_04709_),
    .B(_04710_),
    .C(_04715_),
    .Y(_04716_));
 sky130_fd_sc_hd__nand2_1 _10813_ (.A(_04714_),
    .B(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__inv_2 _10814_ (.A(_04717_),
    .Y(_04718_));
 sky130_fd_sc_hd__nand2_1 _10815_ (.A(_04646_),
    .B(_04718_),
    .Y(_04719_));
 sky130_fd_sc_hd__nand3_1 _10816_ (.A(_04717_),
    .B(_04526_),
    .C(_04645_),
    .Y(_04720_));
 sky130_fd_sc_hd__nand2_1 _10817_ (.A(_04719_),
    .B(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__nand2_1 _10818_ (.A(_04721_),
    .B(_03746_),
    .Y(_04722_));
 sky130_fd_sc_hd__nand2_1 _10819_ (.A(_04600_),
    .B(_04597_),
    .Y(_04723_));
 sky130_fd_sc_hd__nand2_1 _10820_ (.A(_04571_),
    .B(_04568_),
    .Y(_04724_));
 sky130_fd_sc_hd__nor2_1 _10821_ (.A(_03899_),
    .B(_04691_),
    .Y(_04725_));
 sky130_fd_sc_hd__a21oi_1 _10822_ (.A1(_04558_),
    .A2(_04539_),
    .B1(_04557_),
    .Y(_04726_));
 sky130_fd_sc_hd__nor2_1 _10823_ (.A(_04345_),
    .B(_04495_),
    .Y(_04727_));
 sky130_fd_sc_hd__inv_2 _10824_ (.A(_03866_),
    .Y(_04728_));
 sky130_fd_sc_hd__buf_4 _10825_ (.A(_04105_),
    .X(_04729_));
 sky130_fd_sc_hd__nor2_1 _10826_ (.A(_04729_),
    .B(_02416_),
    .Y(_04730_));
 sky130_fd_sc_hd__nand2_1 _10827_ (.A(_04105_),
    .B(\Oset[1][11] ),
    .Y(_04731_));
 sky130_fd_sc_hd__inv_2 _10828_ (.A(_04731_),
    .Y(_04732_));
 sky130_fd_sc_hd__nor2_1 _10829_ (.A(_04105_),
    .B(_02413_),
    .Y(_04733_));
 sky130_fd_sc_hd__a211o_1 _10830_ (.A1(_04729_),
    .A2(\Oset[3][11] ),
    .B1(_04045_),
    .C1(_04733_),
    .X(_04734_));
 sky130_fd_sc_hd__o31ai_4 _10831_ (.A1(_04042_),
    .A2(_04730_),
    .A3(_04732_),
    .B1(_04734_),
    .Y(_04735_));
 sky130_fd_sc_hd__a21oi_1 _10832_ (.A1(_04735_),
    .A2(_03781_),
    .B1(_00585_),
    .Y(_04736_));
 sky130_fd_sc_hd__nor2_1 _10833_ (.A(_04729_),
    .B(_02406_),
    .Y(_04737_));
 sky130_fd_sc_hd__a211o_1 _10834_ (.A1(_04729_),
    .A2(\Qset[3][11] ),
    .B1(_04045_),
    .C1(_04737_),
    .X(_04738_));
 sky130_fd_sc_hd__nor2_1 _10835_ (.A(_04729_),
    .B(_02409_),
    .Y(_04739_));
 sky130_fd_sc_hd__a211o_1 _10836_ (.A1(_04729_),
    .A2(\Qset[1][11] ),
    .B1(_04042_),
    .C1(_04739_),
    .X(_04740_));
 sky130_fd_sc_hd__nand2_2 _10837_ (.A(_04738_),
    .B(_04740_),
    .Y(_04741_));
 sky130_fd_sc_hd__o21ai_1 _10838_ (.A1(_02163_),
    .A2(_04741_),
    .B1(_02872_),
    .Y(_04742_));
 sky130_fd_sc_hd__nand2_1 _10839_ (.A(_04736_),
    .B(_04742_),
    .Y(_04743_));
 sky130_fd_sc_hd__a221oi_4 _10840_ (.A1(_03768_),
    .A2(_04728_),
    .B1(_04743_),
    .B2(_02885_),
    .C1(_00589_),
    .Y(_04744_));
 sky130_fd_sc_hd__nand2_1 _10841_ (.A(_04308_),
    .B(_04744_),
    .Y(_04745_));
 sky130_fd_sc_hd__inv_2 _10842_ (.A(_04744_),
    .Y(_04746_));
 sky130_fd_sc_hd__nand2_1 _10843_ (.A(_04308_),
    .B(_04555_),
    .Y(_04747_));
 sky130_fd_sc_hd__o21ai_1 _10844_ (.A1(_04746_),
    .A2(_04025_),
    .B1(_04747_),
    .Y(_04748_));
 sky130_fd_sc_hd__o21ai_1 _10845_ (.A1(_04556_),
    .A2(_04745_),
    .B1(_04748_),
    .Y(_04749_));
 sky130_fd_sc_hd__xor2_1 _10846_ (.A(_04727_),
    .B(_04749_),
    .X(_04750_));
 sky130_fd_sc_hd__or2_1 _10847_ (.A(_04726_),
    .B(_04750_),
    .X(_04751_));
 sky130_fd_sc_hd__nand2_1 _10848_ (.A(_04750_),
    .B(_04726_),
    .Y(_04752_));
 sky130_fd_sc_hd__nand2_1 _10849_ (.A(_04751_),
    .B(_04752_),
    .Y(_04753_));
 sky130_fd_sc_hd__xor2_1 _10850_ (.A(_04725_),
    .B(_04753_),
    .X(_04754_));
 sky130_fd_sc_hd__a21o_1 _10851_ (.A1(_04561_),
    .A2(_04564_),
    .B1(_04754_),
    .X(_04755_));
 sky130_fd_sc_hd__nand3_1 _10852_ (.A(_04754_),
    .B(_04561_),
    .C(_04564_),
    .Y(_04756_));
 sky130_fd_sc_hd__nand2_2 _10853_ (.A(_04755_),
    .B(_04756_),
    .Y(_04757_));
 sky130_fd_sc_hd__inv_2 _10854_ (.A(_04757_),
    .Y(_04758_));
 sky130_fd_sc_hd__nand2_1 _10855_ (.A(_04724_),
    .B(_04758_),
    .Y(_04759_));
 sky130_fd_sc_hd__nand3_1 _10856_ (.A(_04571_),
    .B(_04568_),
    .C(_04757_),
    .Y(_04760_));
 sky130_fd_sc_hd__nand2_1 _10857_ (.A(_04593_),
    .B(_04589_),
    .Y(_04761_));
 sky130_fd_sc_hd__a21oi_1 _10858_ (.A1(_04584_),
    .A2(_04575_),
    .B1(_04583_),
    .Y(_04762_));
 sky130_fd_sc_hd__nor2_1 _10859_ (.A(_04110_),
    .B(_03685_),
    .Y(_04763_));
 sky130_fd_sc_hd__a21oi_1 _10860_ (.A1(_04580_),
    .A2(_04577_),
    .B1(_04579_),
    .Y(_04764_));
 sky130_fd_sc_hd__nor2_1 _10861_ (.A(_03507_),
    .B(_04050_),
    .Y(_04765_));
 sky130_fd_sc_hd__nand2_1 _10862_ (.A(_04074_),
    .B(_03421_),
    .Y(_04766_));
 sky130_fd_sc_hd__nor2_1 _10863_ (.A(_04766_),
    .B(_04578_),
    .Y(_04767_));
 sky130_fd_sc_hd__nand2_1 _10864_ (.A(_04578_),
    .B(_04766_),
    .Y(_04768_));
 sky130_fd_sc_hd__and2b_1 _10865_ (.A_N(_04767_),
    .B(_04768_),
    .X(_04769_));
 sky130_fd_sc_hd__xnor2_1 _10866_ (.A(_04765_),
    .B(_04769_),
    .Y(_04770_));
 sky130_fd_sc_hd__nor2_1 _10867_ (.A(_04764_),
    .B(_04770_),
    .Y(_04771_));
 sky130_fd_sc_hd__nand2_1 _10868_ (.A(_04770_),
    .B(_04764_),
    .Y(_04772_));
 sky130_fd_sc_hd__and2b_1 _10869_ (.A_N(_04771_),
    .B(_04772_),
    .X(_04773_));
 sky130_fd_sc_hd__xnor2_1 _10870_ (.A(_04763_),
    .B(_04773_),
    .Y(_04774_));
 sky130_fd_sc_hd__xor2_1 _10871_ (.A(_04762_),
    .B(_04774_),
    .X(_04775_));
 sky130_fd_sc_hd__nand2_1 _10872_ (.A(_04761_),
    .B(_04775_),
    .Y(_04776_));
 sky130_fd_sc_hd__nand3b_1 _10873_ (.A_N(_04775_),
    .B(_04593_),
    .C(_04589_),
    .Y(_04777_));
 sky130_fd_sc_hd__nand2_1 _10874_ (.A(_04776_),
    .B(_04777_),
    .Y(_04778_));
 sky130_fd_sc_hd__inv_2 _10875_ (.A(_04778_),
    .Y(_04779_));
 sky130_fd_sc_hd__nand3_1 _10876_ (.A(_04759_),
    .B(_04760_),
    .C(_04779_),
    .Y(_04780_));
 sky130_fd_sc_hd__nand2_1 _10877_ (.A(_04724_),
    .B(_04757_),
    .Y(_04781_));
 sky130_fd_sc_hd__nand3_1 _10878_ (.A(_04571_),
    .B(_04568_),
    .C(_04758_),
    .Y(_04782_));
 sky130_fd_sc_hd__nand3_1 _10879_ (.A(_04781_),
    .B(_04782_),
    .C(_04778_),
    .Y(_04783_));
 sky130_fd_sc_hd__nand2_1 _10880_ (.A(_04780_),
    .B(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__inv_2 _10881_ (.A(_04784_),
    .Y(_04785_));
 sky130_fd_sc_hd__nand2_1 _10882_ (.A(_04723_),
    .B(_04785_),
    .Y(_04786_));
 sky130_fd_sc_hd__nand3_1 _10883_ (.A(_04600_),
    .B(_04784_),
    .C(_04597_),
    .Y(_04787_));
 sky130_fd_sc_hd__nand3_1 _10884_ (.A(_04786_),
    .B(_03048_),
    .C(_04787_),
    .Y(_04788_));
 sky130_fd_sc_hd__a31o_1 _10885_ (.A1(_04759_),
    .A2(_04760_),
    .A3(_03751_),
    .B1(_03745_),
    .X(_04789_));
 sky130_fd_sc_hd__inv_2 _10886_ (.A(_04789_),
    .Y(_04790_));
 sky130_fd_sc_hd__nand2_1 _10887_ (.A(_04788_),
    .B(_04790_),
    .Y(_04791_));
 sky130_fd_sc_hd__nand3_1 _10888_ (.A(_04722_),
    .B(_04791_),
    .C(_00820_),
    .Y(_04792_));
 sky130_fd_sc_hd__nand2_1 _10889_ (.A(_04744_),
    .B(_02096_),
    .Y(_04793_));
 sky130_fd_sc_hd__nand2_1 _10890_ (.A(_04792_),
    .B(_04793_),
    .Y(_04794_));
 sky130_fd_sc_hd__nand2_1 _10891_ (.A(_04794_),
    .B(_02160_),
    .Y(_04795_));
 sky130_fd_sc_hd__nand3_1 _10892_ (.A(_04792_),
    .B(_00831_),
    .C(_04793_),
    .Y(_04796_));
 sky130_fd_sc_hd__a21o_1 _10893_ (.A1(\H[3][11] ),
    .A2(_03793_),
    .B1(_03795_),
    .X(_04797_));
 sky130_fd_sc_hd__a21o_1 _10894_ (.A1(\H[2][11] ),
    .A2(_04415_),
    .B1(_04797_),
    .X(_04798_));
 sky130_fd_sc_hd__nor2_1 _10895_ (.A(_03793_),
    .B(_03861_),
    .Y(_04799_));
 sky130_fd_sc_hd__a211o_1 _10896_ (.A1(\H[1][11] ),
    .A2(_03793_),
    .B1(_03798_),
    .C1(_04799_),
    .X(_04800_));
 sky130_fd_sc_hd__nand2_1 _10897_ (.A(_04414_),
    .B(\Qset[0][11] ),
    .Y(_04801_));
 sky130_fd_sc_hd__nand2_1 _10898_ (.A(\Qset[1][11] ),
    .B(_03792_),
    .Y(_04802_));
 sky130_fd_sc_hd__a21oi_1 _10899_ (.A1(\Qset[3][11] ),
    .A2(_03792_),
    .B1(_03795_),
    .Y(_04803_));
 sky130_fd_sc_hd__nand2_1 _10900_ (.A(_04415_),
    .B(\Qset[2][11] ),
    .Y(_04804_));
 sky130_fd_sc_hd__a32o_1 _10901_ (.A1(_04801_),
    .A2(_04802_),
    .A3(_03795_),
    .B1(_04803_),
    .B2(_04804_),
    .X(_04805_));
 sky130_fd_sc_hd__nand2_1 _10902_ (.A(_04414_),
    .B(\Oset[0][11] ),
    .Y(_04806_));
 sky130_fd_sc_hd__nand2_1 _10903_ (.A(\Oset[1][11] ),
    .B(_03792_),
    .Y(_04807_));
 sky130_fd_sc_hd__a21oi_1 _10904_ (.A1(\Oset[3][11] ),
    .A2(_03792_),
    .B1(_03795_),
    .Y(_04808_));
 sky130_fd_sc_hd__nand2_1 _10905_ (.A(_04414_),
    .B(\Oset[2][11] ),
    .Y(_04809_));
 sky130_fd_sc_hd__a32o_1 _10906_ (.A1(_04806_),
    .A2(_04807_),
    .A3(_03795_),
    .B1(_04808_),
    .B2(_04809_),
    .X(_04810_));
 sky130_fd_sc_hd__mux2_1 _10907_ (.A0(_04805_),
    .A1(_04810_),
    .S(_00621_),
    .X(_04811_));
 sky130_fd_sc_hd__nor2_1 _10908_ (.A(_01538_),
    .B(_04811_),
    .Y(_04812_));
 sky130_fd_sc_hd__a311o_2 _10909_ (.A1(_01538_),
    .A2(_04798_),
    .A3(_04800_),
    .B1(_00556_),
    .C1(_04812_),
    .X(_04813_));
 sky130_fd_sc_hd__o21ai_2 _10910_ (.A1(_00710_),
    .A2(_04690_),
    .B1(_04813_),
    .Y(_04814_));
 sky130_fd_sc_hd__inv_2 _10911_ (.A(_04814_),
    .Y(_04815_));
 sky130_fd_sc_hd__nand3_2 _10912_ (.A(_04795_),
    .B(_04796_),
    .C(_04815_),
    .Y(_04816_));
 sky130_fd_sc_hd__nand2_1 _10913_ (.A(_04794_),
    .B(_00832_),
    .Y(_04817_));
 sky130_fd_sc_hd__nand3_1 _10914_ (.A(_04792_),
    .B(_02160_),
    .C(_04793_),
    .Y(_04818_));
 sky130_fd_sc_hd__nand3_1 _10915_ (.A(_04817_),
    .B(_04818_),
    .C(_04814_),
    .Y(_04819_));
 sky130_fd_sc_hd__nand2_1 _10916_ (.A(_04816_),
    .B(_04819_),
    .Y(_04820_));
 sky130_fd_sc_hd__inv_2 _10917_ (.A(_04633_),
    .Y(_04821_));
 sky130_fd_sc_hd__nand2_1 _10918_ (.A(_04820_),
    .B(_04821_),
    .Y(_04822_));
 sky130_fd_sc_hd__nand3_1 _10919_ (.A(_04816_),
    .B(_04819_),
    .C(_04633_),
    .Y(_04823_));
 sky130_fd_sc_hd__nand2_2 _10920_ (.A(_04822_),
    .B(_04823_),
    .Y(_04824_));
 sky130_fd_sc_hd__nand2_1 _10921_ (.A(_04641_),
    .B(_04636_),
    .Y(_04825_));
 sky130_fd_sc_hd__xor2_2 _10922_ (.A(_04824_),
    .B(_04825_),
    .X(_04826_));
 sky130_fd_sc_hd__clkbuf_4 _10923_ (.A(_00472_),
    .X(_04827_));
 sky130_fd_sc_hd__o21a_1 _10924_ (.A1(\result_reg_add[11] ),
    .A2(_02649_),
    .B1(_04827_),
    .X(_04828_));
 sky130_fd_sc_hd__o21ai_1 _10925_ (.A1(_02654_),
    .A2(_04826_),
    .B1(_04828_),
    .Y(_04829_));
 sky130_fd_sc_hd__inv_2 _10926_ (.A(_04829_),
    .Y(_00255_));
 sky130_fd_sc_hd__buf_6 _10927_ (.A(_00820_),
    .X(_04830_));
 sky130_fd_sc_hd__or2_1 _10928_ (.A(_04283_),
    .B(\H[0][12] ),
    .X(_04831_));
 sky130_fd_sc_hd__buf_6 _10929_ (.A(_04283_),
    .X(_04832_));
 sky130_fd_sc_hd__a21oi_1 _10930_ (.A1(_02446_),
    .A2(_04832_),
    .B1(_03764_),
    .Y(_04833_));
 sky130_fd_sc_hd__mux2_1 _10931_ (.A0(\H[2][12] ),
    .A1(\H[3][12] ),
    .S(_04283_),
    .X(_04834_));
 sky130_fd_sc_hd__clkbuf_4 _10932_ (.A(_03764_),
    .X(_04835_));
 sky130_fd_sc_hd__a22o_1 _10933_ (.A1(_04831_),
    .A2(_04833_),
    .B1(_04834_),
    .B2(_04835_),
    .X(_04836_));
 sky130_fd_sc_hd__nand2_1 _10934_ (.A(_03773_),
    .B(_02436_),
    .Y(_04837_));
 sky130_fd_sc_hd__inv_2 _10935_ (.A(\Oset[3][12] ),
    .Y(_04838_));
 sky130_fd_sc_hd__nand2_1 _10936_ (.A(_04838_),
    .B(_03760_),
    .Y(_04839_));
 sky130_fd_sc_hd__o21a_1 _10937_ (.A1(\Oset[1][12] ),
    .A2(_03773_),
    .B1(_03761_),
    .X(_04840_));
 sky130_fd_sc_hd__nand2_1 _10938_ (.A(_03773_),
    .B(_02439_),
    .Y(_04841_));
 sky130_fd_sc_hd__a32o_1 _10939_ (.A1(_04837_),
    .A2(_04839_),
    .A3(_03764_),
    .B1(_04840_),
    .B2(_04841_),
    .X(_04842_));
 sky130_fd_sc_hd__nor2_1 _10940_ (.A(\Qset[3][12] ),
    .B(_03773_),
    .Y(_04843_));
 sky130_fd_sc_hd__o21ai_1 _10941_ (.A1(_03759_),
    .A2(\Qset[2][12] ),
    .B1(_03345_),
    .Y(_04844_));
 sky130_fd_sc_hd__nor2_1 _10942_ (.A(_03759_),
    .B(\Qset[0][12] ),
    .Y(_04845_));
 sky130_fd_sc_hd__o21ai_1 _10943_ (.A1(\Qset[1][12] ),
    .A2(_03773_),
    .B1(_03004_),
    .Y(_04846_));
 sky130_fd_sc_hd__o22a_1 _10944_ (.A1(_04843_),
    .A2(_04844_),
    .B1(_04845_),
    .B2(_04846_),
    .X(_04847_));
 sky130_fd_sc_hd__and2_1 _10945_ (.A(_04847_),
    .B(_00582_),
    .X(_04848_));
 sky130_fd_sc_hd__a211oi_1 _10946_ (.A1(_02162_),
    .A2(_02435_),
    .B1(_03781_),
    .C1(_04848_),
    .Y(_04849_));
 sky130_fd_sc_hd__a211o_1 _10947_ (.A1(_03781_),
    .A2(_04842_),
    .B1(_00584_),
    .C1(_04849_),
    .X(_04850_));
 sky130_fd_sc_hd__a21oi_1 _10948_ (.A1(_02442_),
    .A2(_00585_),
    .B1(_03768_),
    .Y(_04851_));
 sky130_fd_sc_hd__a22o_1 _10949_ (.A1(_03768_),
    .A2(_04836_),
    .B1(_04850_),
    .B2(_04851_),
    .X(_04852_));
 sky130_fd_sc_hd__nand2_2 _10950_ (.A(_04852_),
    .B(_01553_),
    .Y(_04853_));
 sky130_fd_sc_hd__nand2_8 _10951_ (.A(_04853_),
    .B(_02449_),
    .Y(_04854_));
 sky130_fd_sc_hd__buf_2 _10952_ (.A(_04415_),
    .X(_04855_));
 sky130_fd_sc_hd__buf_2 _10953_ (.A(_04855_),
    .X(_04856_));
 sky130_fd_sc_hd__clkbuf_4 _10954_ (.A(_03793_),
    .X(_04857_));
 sky130_fd_sc_hd__clkbuf_4 _10955_ (.A(_04857_),
    .X(_04858_));
 sky130_fd_sc_hd__clkbuf_4 _10956_ (.A(_03795_),
    .X(_04859_));
 sky130_fd_sc_hd__a21o_1 _10957_ (.A1(\H[3][12] ),
    .A2(_04858_),
    .B1(_04859_),
    .X(_04860_));
 sky130_fd_sc_hd__a21o_1 _10958_ (.A1(\H[2][12] ),
    .A2(_04856_),
    .B1(_04860_),
    .X(_04861_));
 sky130_fd_sc_hd__clkbuf_4 _10959_ (.A(_03798_),
    .X(_04862_));
 sky130_fd_sc_hd__a21oi_1 _10960_ (.A1(_04856_),
    .A2(\H[0][12] ),
    .B1(_04862_),
    .Y(_04863_));
 sky130_fd_sc_hd__o21ai_1 _10961_ (.A1(_02446_),
    .A2(_04856_),
    .B1(_04863_),
    .Y(_04864_));
 sky130_fd_sc_hd__nand2_1 _10962_ (.A(\Oset[1][12] ),
    .B(_04858_),
    .Y(_04865_));
 sky130_fd_sc_hd__a21oi_1 _10963_ (.A1(_04856_),
    .A2(\Oset[0][12] ),
    .B1(_04862_),
    .Y(_04866_));
 sky130_fd_sc_hd__mux2_1 _10964_ (.A0(_02436_),
    .A1(_04838_),
    .S(_04858_),
    .X(_04867_));
 sky130_fd_sc_hd__a221o_1 _10965_ (.A1(_04865_),
    .A2(_04866_),
    .B1(_04867_),
    .B2(_04862_),
    .C1(_00647_),
    .X(_04868_));
 sky130_fd_sc_hd__a21oi_1 _10966_ (.A1(\Qset[3][12] ),
    .A2(_04858_),
    .B1(_04859_),
    .Y(_04869_));
 sky130_fd_sc_hd__nand2_1 _10967_ (.A(_04856_),
    .B(\Qset[2][12] ),
    .Y(_04870_));
 sky130_fd_sc_hd__a21oi_1 _10968_ (.A1(_04856_),
    .A2(\Qset[0][12] ),
    .B1(_04862_),
    .Y(_04871_));
 sky130_fd_sc_hd__nand2_1 _10969_ (.A(\Qset[1][12] ),
    .B(_04858_),
    .Y(_04872_));
 sky130_fd_sc_hd__a221o_1 _10970_ (.A1(_04869_),
    .A2(_04870_),
    .B1(_04871_),
    .B2(_04872_),
    .C1(_00621_),
    .X(_04873_));
 sky130_fd_sc_hd__a21oi_1 _10971_ (.A1(_04868_),
    .A2(_04873_),
    .B1(_01538_),
    .Y(_04874_));
 sky130_fd_sc_hd__a311o_2 _10972_ (.A1(_01538_),
    .A2(_04861_),
    .A3(_04864_),
    .B1(_02096_),
    .C1(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__o21a_1 _10973_ (.A1(_04830_),
    .A2(_04854_),
    .B1(_04875_),
    .X(_04876_));
 sky130_fd_sc_hd__clkinvlp_2 _10974_ (.A(_04816_),
    .Y(_04877_));
 sky130_fd_sc_hd__nand3_1 _10975_ (.A(_04825_),
    .B(_04877_),
    .C(_04824_),
    .Y(_04878_));
 sky130_fd_sc_hd__nand2_1 _10976_ (.A(_04878_),
    .B(_03274_),
    .Y(_04879_));
 sky130_fd_sc_hd__inv_2 _10977_ (.A(_04879_),
    .Y(_04880_));
 sky130_fd_sc_hd__buf_4 _10978_ (.A(_04729_),
    .X(_04881_));
 sky130_fd_sc_hd__nand2_1 _10979_ (.A(_04881_),
    .B(\Oset[1][12] ),
    .Y(_04882_));
 sky130_fd_sc_hd__a21oi_1 _10980_ (.A1(_03152_),
    .A2(\Oset[0][12] ),
    .B1(_04042_),
    .Y(_04883_));
 sky130_fd_sc_hd__nor2_1 _10981_ (.A(_04881_),
    .B(_02436_),
    .Y(_04884_));
 sky130_fd_sc_hd__a21o_1 _10982_ (.A1(_04729_),
    .A2(\Oset[3][12] ),
    .B1(_04045_),
    .X(_04885_));
 sky130_fd_sc_hd__o2bb2a_1 _10983_ (.A1_N(_04882_),
    .A2_N(_04883_),
    .B1(_04884_),
    .B2(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__o21a_1 _10984_ (.A1(_03770_),
    .A2(_04886_),
    .B1(_01156_),
    .X(_04887_));
 sky130_fd_sc_hd__mux2_1 _10985_ (.A0(\Qset[2][12] ),
    .A1(\Qset[3][12] ),
    .S(_04729_),
    .X(_04888_));
 sky130_fd_sc_hd__nor2_1 _10986_ (.A(_04881_),
    .B(_02432_),
    .Y(_04889_));
 sky130_fd_sc_hd__a211o_1 _10987_ (.A1(_04881_),
    .A2(\Qset[1][12] ),
    .B1(_04042_),
    .C1(_04889_),
    .X(_04890_));
 sky130_fd_sc_hd__o21ai_4 _10988_ (.A1(_04045_),
    .A2(_04888_),
    .B1(_04890_),
    .Y(_04891_));
 sky130_fd_sc_hd__o21ai_1 _10989_ (.A1(_02163_),
    .A2(_04891_),
    .B1(_02542_),
    .Y(_04892_));
 sky130_fd_sc_hd__a221o_2 _10990_ (.A1(_00498_),
    .A2(_00585_),
    .B1(_04887_),
    .B2(_04892_),
    .C1(_03768_),
    .X(_04893_));
 sky130_fd_sc_hd__nand2_1 _10991_ (.A(_04108_),
    .B(_03745_),
    .Y(_04894_));
 sky130_fd_sc_hd__nand2_2 _10992_ (.A(_04893_),
    .B(_04894_),
    .Y(_04895_));
 sky130_fd_sc_hd__inv_4 _10993_ (.A(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__nand2_1 _10994_ (.A(_04786_),
    .B(_04780_),
    .Y(_04897_));
 sky130_fd_sc_hd__a21oi_1 _10995_ (.A1(_04772_),
    .A2(_04763_),
    .B1(_04771_),
    .Y(_04898_));
 sky130_fd_sc_hd__nand2_2 _10996_ (.A(_04896_),
    .B(_03079_),
    .Y(_04899_));
 sky130_fd_sc_hd__a21oi_1 _10997_ (.A1(_04768_),
    .A2(_04765_),
    .B1(_04767_),
    .Y(_04900_));
 sky130_fd_sc_hd__nand2_1 _10998_ (.A(_04096_),
    .B(_03506_),
    .Y(_04901_));
 sky130_fd_sc_hd__a22o_1 _10999_ (.A1(_04074_),
    .A2(_03506_),
    .B1(_04096_),
    .B2(_03421_),
    .X(_04902_));
 sky130_fd_sc_hd__o21ai_1 _11000_ (.A1(_04766_),
    .A2(_04901_),
    .B1(_04902_),
    .Y(_04903_));
 sky130_fd_sc_hd__or3_1 _11001_ (.A(_03685_),
    .B(_04050_),
    .C(_04903_),
    .X(_04904_));
 sky130_fd_sc_hd__o21ai_1 _11002_ (.A1(_03685_),
    .A2(_04050_),
    .B1(_04903_),
    .Y(_04905_));
 sky130_fd_sc_hd__nand2_1 _11003_ (.A(_04904_),
    .B(_04905_),
    .Y(_04906_));
 sky130_fd_sc_hd__or2_1 _11004_ (.A(_04900_),
    .B(_04906_),
    .X(_04907_));
 sky130_fd_sc_hd__nand2_1 _11005_ (.A(_04906_),
    .B(_04900_),
    .Y(_04908_));
 sky130_fd_sc_hd__nand2_1 _11006_ (.A(_04907_),
    .B(_04908_),
    .Y(_04909_));
 sky130_fd_sc_hd__or3_1 _11007_ (.A(_04025_),
    .B(_04899_),
    .C(_04909_),
    .X(_04910_));
 sky130_fd_sc_hd__o21ai_1 _11008_ (.A1(_04025_),
    .A2(_04899_),
    .B1(_04909_),
    .Y(_04911_));
 sky130_fd_sc_hd__nand2_1 _11009_ (.A(_04910_),
    .B(_04911_),
    .Y(_04912_));
 sky130_fd_sc_hd__or2_1 _11010_ (.A(_04898_),
    .B(_04912_),
    .X(_04913_));
 sky130_fd_sc_hd__nand2_1 _11011_ (.A(_04912_),
    .B(_04898_),
    .Y(_04914_));
 sky130_fd_sc_hd__nand2_1 _11012_ (.A(_04913_),
    .B(_04914_),
    .Y(_04915_));
 sky130_fd_sc_hd__inv_2 _11013_ (.A(_04915_),
    .Y(_04916_));
 sky130_fd_sc_hd__o21ai_1 _11014_ (.A1(_04762_),
    .A2(_04774_),
    .B1(_04776_),
    .Y(_04917_));
 sky130_fd_sc_hd__or2_1 _11015_ (.A(_04916_),
    .B(_04917_),
    .X(_04918_));
 sky130_fd_sc_hd__nand2_1 _11016_ (.A(_04917_),
    .B(_04916_),
    .Y(_04919_));
 sky130_fd_sc_hd__nand2_1 _11017_ (.A(_04918_),
    .B(_04919_),
    .Y(_04920_));
 sky130_fd_sc_hd__or2_1 _11018_ (.A(_04757_),
    .B(_04571_),
    .X(_04921_));
 sky130_fd_sc_hd__o21a_1 _11019_ (.A1(_04568_),
    .A2(_04757_),
    .B1(_04755_),
    .X(_04922_));
 sky130_fd_sc_hd__o31a_1 _11020_ (.A1(_03899_),
    .A2(_04691_),
    .A3(_04753_),
    .B1(_04751_),
    .X(_04923_));
 sky130_fd_sc_hd__clkinv_4 _11021_ (.A(_04854_),
    .Y(_04924_));
 sky130_fd_sc_hd__nor2_1 _11022_ (.A(_03233_),
    .B(_03899_),
    .Y(_04925_));
 sky130_fd_sc_hd__inv_2 _11023_ (.A(_04925_),
    .Y(_04926_));
 sky130_fd_sc_hd__o2bb2a_1 _11024_ (.A1_N(_04748_),
    .A2_N(_04727_),
    .B1(_04556_),
    .B2(_04745_),
    .X(_04927_));
 sky130_fd_sc_hd__nand2_1 _11025_ (.A(_04690_),
    .B(_03859_),
    .Y(_04928_));
 sky130_fd_sc_hd__nand2_1 _11026_ (.A(_04494_),
    .B(_04744_),
    .Y(_04929_));
 sky130_fd_sc_hd__o21ai_1 _11027_ (.A1(_04607_),
    .A2(_04495_),
    .B1(_04745_),
    .Y(_04930_));
 sky130_fd_sc_hd__o21ai_1 _11028_ (.A1(_04747_),
    .A2(_04929_),
    .B1(_04930_),
    .Y(_04931_));
 sky130_fd_sc_hd__or2_1 _11029_ (.A(_04928_),
    .B(_04931_),
    .X(_04932_));
 sky130_fd_sc_hd__nand2_1 _11030_ (.A(_04931_),
    .B(_04928_),
    .Y(_04933_));
 sky130_fd_sc_hd__nand2_1 _11031_ (.A(_04932_),
    .B(_04933_),
    .Y(_04934_));
 sky130_fd_sc_hd__or2_1 _11032_ (.A(_04927_),
    .B(_04934_),
    .X(_04935_));
 sky130_fd_sc_hd__nand2_1 _11033_ (.A(_04934_),
    .B(_04927_),
    .Y(_04936_));
 sky130_fd_sc_hd__nand2_1 _11034_ (.A(_04935_),
    .B(_04936_),
    .Y(_04937_));
 sky130_fd_sc_hd__or3_1 _11035_ (.A(_04924_),
    .B(_04926_),
    .C(_04937_),
    .X(_04938_));
 sky130_fd_sc_hd__o21ai_1 _11036_ (.A1(_04924_),
    .A2(_04926_),
    .B1(_04937_),
    .Y(_04939_));
 sky130_fd_sc_hd__nand2_1 _11037_ (.A(_04938_),
    .B(_04939_),
    .Y(_04940_));
 sky130_fd_sc_hd__or2_1 _11038_ (.A(_04923_),
    .B(_04940_),
    .X(_04941_));
 sky130_fd_sc_hd__nand2_1 _11039_ (.A(_04940_),
    .B(_04923_),
    .Y(_04942_));
 sky130_fd_sc_hd__nand2_1 _11040_ (.A(_04941_),
    .B(_04942_),
    .Y(_04943_));
 sky130_fd_sc_hd__a21o_1 _11041_ (.A1(_04921_),
    .A2(_04922_),
    .B1(_04943_),
    .X(_04944_));
 sky130_fd_sc_hd__nand3_1 _11042_ (.A(_04921_),
    .B(_04922_),
    .C(_04943_),
    .Y(_04945_));
 sky130_fd_sc_hd__nand2_1 _11043_ (.A(_04944_),
    .B(_04945_),
    .Y(_04946_));
 sky130_fd_sc_hd__or2_1 _11044_ (.A(_04920_),
    .B(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__nand2_1 _11045_ (.A(_04946_),
    .B(_04920_),
    .Y(_04948_));
 sky130_fd_sc_hd__nand2_1 _11046_ (.A(_04947_),
    .B(_04948_),
    .Y(_04949_));
 sky130_fd_sc_hd__inv_2 _11047_ (.A(_04949_),
    .Y(_04950_));
 sky130_fd_sc_hd__or2_1 _11048_ (.A(_04897_),
    .B(_04950_),
    .X(_04951_));
 sky130_fd_sc_hd__nand2_1 _11049_ (.A(_04950_),
    .B(_04897_),
    .Y(_04952_));
 sky130_fd_sc_hd__a21o_1 _11050_ (.A1(_04951_),
    .A2(_04952_),
    .B1(_03751_),
    .X(_04953_));
 sky130_fd_sc_hd__nand2_1 _11051_ (.A(_03652_),
    .B(_04096_),
    .Y(_04954_));
 sky130_fd_sc_hd__inv_2 _11052_ (.A(_04073_),
    .Y(_04955_));
 sky130_fd_sc_hd__nand2_1 _11053_ (.A(_04955_),
    .B(_03079_),
    .Y(_04956_));
 sky130_fd_sc_hd__inv_2 _11054_ (.A(_04956_),
    .Y(_04957_));
 sky130_fd_sc_hd__nand2_1 _11055_ (.A(_03790_),
    .B(_04957_),
    .Y(_04958_));
 sky130_fd_sc_hd__nor2_1 _11056_ (.A(_04954_),
    .B(_04958_),
    .Y(_04959_));
 sky130_fd_sc_hd__mux2_1 _11057_ (.A0(\Qset[2][13] ),
    .A1(\Qset[3][13] ),
    .S(_04729_),
    .X(_04960_));
 sky130_fd_sc_hd__nor2_1 _11058_ (.A(_04881_),
    .B(_02455_),
    .Y(_04961_));
 sky130_fd_sc_hd__a211o_1 _11059_ (.A1(_04881_),
    .A2(\Qset[1][13] ),
    .B1(_04042_),
    .C1(_04961_),
    .X(_04962_));
 sky130_fd_sc_hd__o21ai_4 _11060_ (.A1(_04045_),
    .A2(_04960_),
    .B1(_04962_),
    .Y(_04963_));
 sky130_fd_sc_hd__o21ai_1 _11061_ (.A1(_02163_),
    .A2(_04963_),
    .B1(_02713_),
    .Y(_04964_));
 sky130_fd_sc_hd__nor2_1 _11062_ (.A(_04881_),
    .B(_02463_),
    .Y(_04965_));
 sky130_fd_sc_hd__a211o_1 _11063_ (.A1(_04881_),
    .A2(\Oset[1][13] ),
    .B1(_04042_),
    .C1(_04965_),
    .X(_04966_));
 sky130_fd_sc_hd__nor2_1 _11064_ (.A(_04881_),
    .B(_02460_),
    .Y(_04967_));
 sky130_fd_sc_hd__a211o_1 _11065_ (.A1(_04881_),
    .A2(\Oset[3][13] ),
    .B1(_04045_),
    .C1(_04967_),
    .X(_04968_));
 sky130_fd_sc_hd__nand2_2 _11066_ (.A(_04966_),
    .B(_04968_),
    .Y(_04969_));
 sky130_fd_sc_hd__nand2_1 _11067_ (.A(_04969_),
    .B(_03781_),
    .Y(_04970_));
 sky130_fd_sc_hd__a31o_1 _11068_ (.A1(_04964_),
    .A2(_01156_),
    .A3(_04970_),
    .B1(_03132_),
    .X(_04971_));
 sky130_fd_sc_hd__nand2_1 _11069_ (.A(_04048_),
    .B(_03745_),
    .Y(_04972_));
 sky130_fd_sc_hd__nand2_1 _11070_ (.A(_04971_),
    .B(_04972_),
    .Y(_04973_));
 sky130_fd_sc_hd__inv_2 _11071_ (.A(_04973_),
    .Y(_04974_));
 sky130_fd_sc_hd__nand2_2 _11072_ (.A(_04974_),
    .B(_03079_),
    .Y(_04975_));
 sky130_fd_sc_hd__nand2_1 _11073_ (.A(_04958_),
    .B(_04954_),
    .Y(_04976_));
 sky130_fd_sc_hd__nand2b_1 _11074_ (.A_N(_04959_),
    .B(_04976_),
    .Y(_04977_));
 sky130_fd_sc_hd__or3_1 _11075_ (.A(_04309_),
    .B(_04975_),
    .C(_04977_),
    .X(_04978_));
 sky130_fd_sc_hd__and2b_1 _11076_ (.A_N(_04959_),
    .B(_04978_),
    .X(_04979_));
 sky130_fd_sc_hd__inv_2 _11077_ (.A(_04095_),
    .Y(_04980_));
 sky130_fd_sc_hd__nand2_1 _11078_ (.A(_04980_),
    .B(_03079_),
    .Y(_04981_));
 sky130_fd_sc_hd__inv_2 _11079_ (.A(_04981_),
    .Y(_04982_));
 sky130_fd_sc_hd__nand2_1 _11080_ (.A(_04308_),
    .B(_04982_),
    .Y(_04983_));
 sky130_fd_sc_hd__a22o_1 _11081_ (.A1(_04308_),
    .A2(_04957_),
    .B1(_03790_),
    .B2(_04982_),
    .X(_04984_));
 sky130_fd_sc_hd__o21ai_1 _11082_ (.A1(_04958_),
    .A2(_04983_),
    .B1(_04984_),
    .Y(_04985_));
 sky130_fd_sc_hd__or3_1 _11083_ (.A(_04495_),
    .B(_04975_),
    .C(_04985_),
    .X(_04986_));
 sky130_fd_sc_hd__o21ai_1 _11084_ (.A1(_04495_),
    .A2(_04975_),
    .B1(_04985_),
    .Y(_04987_));
 sky130_fd_sc_hd__nand2_1 _11085_ (.A(_04986_),
    .B(_04987_),
    .Y(_04988_));
 sky130_fd_sc_hd__or2_1 _11086_ (.A(_04979_),
    .B(_04988_),
    .X(_04989_));
 sky130_fd_sc_hd__nand2_1 _11087_ (.A(_04988_),
    .B(_04979_),
    .Y(_04990_));
 sky130_fd_sc_hd__nand2_1 _11088_ (.A(_04989_),
    .B(_04990_),
    .Y(_04991_));
 sky130_fd_sc_hd__or3_1 _11089_ (.A(_04691_),
    .B(_04899_),
    .C(_04991_),
    .X(_04992_));
 sky130_fd_sc_hd__and2_1 _11090_ (.A(_04992_),
    .B(_04989_),
    .X(_04993_));
 sky130_fd_sc_hd__nor2_1 _11091_ (.A(_04975_),
    .B(_04691_),
    .Y(_04994_));
 sky130_fd_sc_hd__nand2_1 _11092_ (.A(_04494_),
    .B(_04957_),
    .Y(_04995_));
 sky130_fd_sc_hd__nor2_1 _11093_ (.A(_04983_),
    .B(_04995_),
    .Y(_04996_));
 sky130_fd_sc_hd__nand2_1 _11094_ (.A(_04995_),
    .B(_04983_),
    .Y(_04997_));
 sky130_fd_sc_hd__and2b_1 _11095_ (.A_N(_04996_),
    .B(_04997_),
    .X(_04998_));
 sky130_fd_sc_hd__xnor2_1 _11096_ (.A(_04994_),
    .B(_04998_),
    .Y(_04999_));
 sky130_fd_sc_hd__o21a_1 _11097_ (.A1(_04958_),
    .A2(_04983_),
    .B1(_04986_),
    .X(_05000_));
 sky130_fd_sc_hd__nor2_1 _11098_ (.A(_04999_),
    .B(_05000_),
    .Y(_05001_));
 sky130_fd_sc_hd__nand2_1 _11099_ (.A(_05000_),
    .B(_04999_),
    .Y(_05002_));
 sky130_fd_sc_hd__or2b_1 _11100_ (.A(_05001_),
    .B_N(_05002_),
    .X(_05003_));
 sky130_fd_sc_hd__or3_1 _11101_ (.A(_04895_),
    .B(_04924_),
    .C(_05003_),
    .X(_05004_));
 sky130_fd_sc_hd__o21ai_1 _11102_ (.A1(_04895_),
    .A2(_04924_),
    .B1(_05003_),
    .Y(_05005_));
 sky130_fd_sc_hd__nand2_1 _11103_ (.A(_05004_),
    .B(_05005_),
    .Y(_05006_));
 sky130_fd_sc_hd__or2_1 _11104_ (.A(_04993_),
    .B(_05006_),
    .X(_05007_));
 sky130_fd_sc_hd__nand2_1 _11105_ (.A(_05006_),
    .B(_04993_),
    .Y(_05008_));
 sky130_fd_sc_hd__and2_1 _11106_ (.A(_05007_),
    .B(_05008_),
    .X(_05009_));
 sky130_fd_sc_hd__nand2_1 _11107_ (.A(_04919_),
    .B(_04913_),
    .Y(_05010_));
 sky130_fd_sc_hd__nor2_1 _11108_ (.A(_04309_),
    .B(_04899_),
    .Y(_05011_));
 sky130_fd_sc_hd__nor2_1 _11109_ (.A(_04975_),
    .B(_04025_),
    .Y(_05012_));
 sky130_fd_sc_hd__nand2_1 _11110_ (.A(_04074_),
    .B(_03506_),
    .Y(_05013_));
 sky130_fd_sc_hd__a21bo_1 _11111_ (.A1(_03652_),
    .A2(_04074_),
    .B1_N(_04901_),
    .X(_05014_));
 sky130_fd_sc_hd__o21ai_1 _11112_ (.A1(_05013_),
    .A2(_04954_),
    .B1(_05014_),
    .Y(_05015_));
 sky130_fd_sc_hd__xor2_1 _11113_ (.A(_05012_),
    .B(_05015_),
    .X(_05016_));
 sky130_fd_sc_hd__o21a_1 _11114_ (.A1(_04766_),
    .A2(_04901_),
    .B1(_04904_),
    .X(_05017_));
 sky130_fd_sc_hd__or2_1 _11115_ (.A(_05016_),
    .B(_05017_),
    .X(_05018_));
 sky130_fd_sc_hd__nand2_1 _11116_ (.A(_05017_),
    .B(_05016_),
    .Y(_05019_));
 sky130_fd_sc_hd__nand2_1 _11117_ (.A(_05018_),
    .B(_05019_),
    .Y(_05020_));
 sky130_fd_sc_hd__xor2_1 _11118_ (.A(_05011_),
    .B(_05020_),
    .X(_05021_));
 sky130_fd_sc_hd__and2_1 _11119_ (.A(_04910_),
    .B(_04907_),
    .X(_05022_));
 sky130_fd_sc_hd__nor2_1 _11120_ (.A(_05021_),
    .B(_05022_),
    .Y(_05023_));
 sky130_fd_sc_hd__inv_2 _11121_ (.A(_05023_),
    .Y(_05024_));
 sky130_fd_sc_hd__nand2_1 _11122_ (.A(_05022_),
    .B(_05021_),
    .Y(_05025_));
 sky130_fd_sc_hd__and2_1 _11123_ (.A(_05024_),
    .B(_05025_),
    .X(_05026_));
 sky130_fd_sc_hd__nand2_1 _11124_ (.A(_05010_),
    .B(_05026_),
    .Y(_05027_));
 sky130_fd_sc_hd__nand2_1 _11125_ (.A(_05027_),
    .B(_05024_),
    .Y(_05028_));
 sky130_fd_sc_hd__nor2_1 _11126_ (.A(_04495_),
    .B(_04899_),
    .Y(_05029_));
 sky130_fd_sc_hd__o2bb2a_1 _11127_ (.A1_N(_05014_),
    .A2_N(_05012_),
    .B1(_05013_),
    .B2(_04954_),
    .X(_05030_));
 sky130_fd_sc_hd__o21ai_1 _11128_ (.A1(_04309_),
    .A2(_04975_),
    .B1(_04977_),
    .Y(_05031_));
 sky130_fd_sc_hd__nand2_1 _11129_ (.A(_04978_),
    .B(_05031_),
    .Y(_05032_));
 sky130_fd_sc_hd__or2_1 _11130_ (.A(_05030_),
    .B(_05032_),
    .X(_05033_));
 sky130_fd_sc_hd__nand2_1 _11131_ (.A(_05032_),
    .B(_05030_),
    .Y(_05034_));
 sky130_fd_sc_hd__nand2_1 _11132_ (.A(_05033_),
    .B(_05034_),
    .Y(_05035_));
 sky130_fd_sc_hd__xor2_1 _11133_ (.A(_05029_),
    .B(_05035_),
    .X(_05036_));
 sky130_fd_sc_hd__o31a_1 _11134_ (.A1(_04309_),
    .A2(_04899_),
    .A3(_05020_),
    .B1(_05018_),
    .X(_05037_));
 sky130_fd_sc_hd__or2_1 _11135_ (.A(_05036_),
    .B(_05037_),
    .X(_05038_));
 sky130_fd_sc_hd__nand2_1 _11136_ (.A(_05037_),
    .B(_05036_),
    .Y(_05039_));
 sky130_fd_sc_hd__nand2_1 _11137_ (.A(_05038_),
    .B(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__inv_2 _11138_ (.A(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__nand2_1 _11139_ (.A(_05028_),
    .B(_05041_),
    .Y(_05042_));
 sky130_fd_sc_hd__nand2_1 _11140_ (.A(_05042_),
    .B(_05038_),
    .Y(_05043_));
 sky130_fd_sc_hd__a21bo_1 _11141_ (.A1(_05029_),
    .A2(_05034_),
    .B1_N(_05033_),
    .X(_05044_));
 sky130_fd_sc_hd__o21ai_1 _11142_ (.A1(_04691_),
    .A2(_04899_),
    .B1(_04991_),
    .Y(_05045_));
 sky130_fd_sc_hd__nand2_1 _11143_ (.A(_04992_),
    .B(_05045_),
    .Y(_05046_));
 sky130_fd_sc_hd__xnor2_1 _11144_ (.A(_05044_),
    .B(_05046_),
    .Y(_05047_));
 sky130_fd_sc_hd__nand2_1 _11145_ (.A(_05043_),
    .B(_05047_),
    .Y(_05048_));
 sky130_fd_sc_hd__or2b_1 _11146_ (.A(_05046_),
    .B_N(_05044_),
    .X(_05049_));
 sky130_fd_sc_hd__nand2_1 _11147_ (.A(_05048_),
    .B(_05049_),
    .Y(_05050_));
 sky130_fd_sc_hd__or2_1 _11148_ (.A(_05009_),
    .B(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__nand2_1 _11149_ (.A(_05050_),
    .B(_05009_),
    .Y(_05052_));
 sky130_fd_sc_hd__a21o_1 _11150_ (.A1(_05051_),
    .A2(_05052_),
    .B1(_03048_),
    .X(_05053_));
 sky130_fd_sc_hd__nand3_1 _11151_ (.A(_04953_),
    .B(_04196_),
    .C(_05053_),
    .Y(_05054_));
 sky130_fd_sc_hd__nand2_1 _11152_ (.A(_04719_),
    .B(_04716_),
    .Y(_05055_));
 sky130_fd_sc_hd__inv_2 _11153_ (.A(_04176_),
    .Y(_05056_));
 sky130_fd_sc_hd__nand2_1 _11154_ (.A(_04175_),
    .B(_04147_),
    .Y(_05057_));
 sky130_fd_sc_hd__nand2_1 _11155_ (.A(_05056_),
    .B(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__inv_2 _11156_ (.A(_05058_),
    .Y(_05059_));
 sky130_fd_sc_hd__nand2_1 _11157_ (.A(_04709_),
    .B(_04702_),
    .Y(_05060_));
 sky130_fd_sc_hd__nand2_1 _11158_ (.A(_03701_),
    .B(_03699_),
    .Y(_05061_));
 sky130_fd_sc_hd__o31a_1 _11159_ (.A1(_03206_),
    .A2(_03685_),
    .A3(_03697_),
    .B1(_03695_),
    .X(_05062_));
 sky130_fd_sc_hd__nand2_1 _11160_ (.A(_03790_),
    .B(_03745_),
    .Y(_05063_));
 sky130_fd_sc_hd__nand2_1 _11161_ (.A(_03652_),
    .B(_03145_),
    .Y(_05064_));
 sky130_fd_sc_hd__nand2_1 _11162_ (.A(_03505_),
    .B(_03076_),
    .Y(_05065_));
 sky130_fd_sc_hd__or2_1 _11163_ (.A(_03690_),
    .B(_05065_),
    .X(_05066_));
 sky130_fd_sc_hd__nand2_1 _11164_ (.A(_03506_),
    .B(_03110_),
    .Y(_05067_));
 sky130_fd_sc_hd__nand2_1 _11165_ (.A(_05067_),
    .B(_03688_),
    .Y(_05068_));
 sky130_fd_sc_hd__nand2_1 _11166_ (.A(_05066_),
    .B(_05068_),
    .Y(_05069_));
 sky130_fd_sc_hd__or2_1 _11167_ (.A(_05064_),
    .B(_05069_),
    .X(_05070_));
 sky130_fd_sc_hd__nand2_1 _11168_ (.A(_05069_),
    .B(_05064_),
    .Y(_05071_));
 sky130_fd_sc_hd__nand2_1 _11169_ (.A(_05070_),
    .B(_05071_),
    .Y(_05072_));
 sky130_fd_sc_hd__o31a_1 _11170_ (.A1(_03383_),
    .A2(_03507_),
    .A3(_03692_),
    .B1(_03689_),
    .X(_05073_));
 sky130_fd_sc_hd__or2_1 _11171_ (.A(_05072_),
    .B(_05073_),
    .X(_05074_));
 sky130_fd_sc_hd__nand2_1 _11172_ (.A(_05073_),
    .B(_05072_),
    .Y(_05075_));
 sky130_fd_sc_hd__nand2_1 _11173_ (.A(_05074_),
    .B(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__or3_1 _11174_ (.A(_03206_),
    .B(_05063_),
    .C(_05076_),
    .X(_05077_));
 sky130_fd_sc_hd__nor2_1 _11175_ (.A(_03897_),
    .B(_03206_),
    .Y(_05078_));
 sky130_fd_sc_hd__inv_2 _11176_ (.A(_05078_),
    .Y(_05079_));
 sky130_fd_sc_hd__o21ai_1 _11177_ (.A1(_04025_),
    .A2(_05079_),
    .B1(_05076_),
    .Y(_05080_));
 sky130_fd_sc_hd__nand2_1 _11178_ (.A(_05077_),
    .B(_05080_),
    .Y(_05081_));
 sky130_fd_sc_hd__nor2_1 _11179_ (.A(_05062_),
    .B(_05081_),
    .Y(_05082_));
 sky130_fd_sc_hd__inv_2 _11180_ (.A(_05082_),
    .Y(_05083_));
 sky130_fd_sc_hd__nand2_1 _11181_ (.A(_05081_),
    .B(_05062_),
    .Y(_05084_));
 sky130_fd_sc_hd__and2_1 _11182_ (.A(_05083_),
    .B(_05084_),
    .X(_05085_));
 sky130_fd_sc_hd__or2_1 _11183_ (.A(_05061_),
    .B(_05085_),
    .X(_05086_));
 sky130_fd_sc_hd__nand2_1 _11184_ (.A(_05085_),
    .B(_05061_),
    .Y(_05087_));
 sky130_fd_sc_hd__nand2_1 _11185_ (.A(_05086_),
    .B(_05087_),
    .Y(_05088_));
 sky130_fd_sc_hd__o21a_1 _11186_ (.A1(_04663_),
    .A2(_04660_),
    .B1(_04693_),
    .X(_05089_));
 sky130_fd_sc_hd__nor2_1 _11187_ (.A(_04281_),
    .B(_04924_),
    .Y(_05090_));
 sky130_fd_sc_hd__a21oi_1 _11188_ (.A1(_04658_),
    .A2(_04654_),
    .B1(_04653_),
    .Y(_05091_));
 sky130_fd_sc_hd__nor2_1 _11189_ (.A(_04458_),
    .B(_04691_),
    .Y(_05092_));
 sky130_fd_sc_hd__nand2_1 _11190_ (.A(_04494_),
    .B(_04651_),
    .Y(_05093_));
 sky130_fd_sc_hd__nand2_1 _11191_ (.A(_04494_),
    .B(_04460_),
    .Y(_05094_));
 sky130_fd_sc_hd__nand2_1 _11192_ (.A(_04308_),
    .B(_04651_),
    .Y(_05095_));
 sky130_fd_sc_hd__nand2_1 _11193_ (.A(_05094_),
    .B(_05095_),
    .Y(_05096_));
 sky130_fd_sc_hd__o21a_1 _11194_ (.A1(_04650_),
    .A2(_05093_),
    .B1(_05096_),
    .X(_05097_));
 sky130_fd_sc_hd__or2_1 _11195_ (.A(_05092_),
    .B(_05097_),
    .X(_05098_));
 sky130_fd_sc_hd__nand2_1 _11196_ (.A(_05097_),
    .B(_05092_),
    .Y(_05099_));
 sky130_fd_sc_hd__nand2_1 _11197_ (.A(_05098_),
    .B(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__xor2_1 _11198_ (.A(_05091_),
    .B(_05100_),
    .X(_05101_));
 sky130_fd_sc_hd__xnor2_1 _11199_ (.A(_05090_),
    .B(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__xor2_1 _11200_ (.A(_05089_),
    .B(_05102_),
    .X(_05103_));
 sky130_fd_sc_hd__o211ai_2 _11201_ (.A1(_04696_),
    .A2(_04695_),
    .B1(_04703_),
    .C1(_04704_),
    .Y(_05104_));
 sky130_fd_sc_hd__xnor2_1 _11202_ (.A(_05103_),
    .B(_05104_),
    .Y(_05105_));
 sky130_fd_sc_hd__xnor2_1 _11203_ (.A(_05088_),
    .B(_05105_),
    .Y(_05106_));
 sky130_fd_sc_hd__inv_2 _11204_ (.A(_05106_),
    .Y(_05107_));
 sky130_fd_sc_hd__or2_1 _11205_ (.A(_05060_),
    .B(_05107_),
    .X(_05108_));
 sky130_fd_sc_hd__nand2_1 _11206_ (.A(_05107_),
    .B(_05060_),
    .Y(_05109_));
 sky130_fd_sc_hd__nand2_1 _11207_ (.A(_05108_),
    .B(_05109_),
    .Y(_05110_));
 sky130_fd_sc_hd__xor2_1 _11208_ (.A(_05059_),
    .B(_05110_),
    .X(_05111_));
 sky130_fd_sc_hd__inv_2 _11209_ (.A(_05111_),
    .Y(_05112_));
 sky130_fd_sc_hd__or2_1 _11210_ (.A(_05055_),
    .B(_05112_),
    .X(_05113_));
 sky130_fd_sc_hd__nand2_1 _11211_ (.A(_05112_),
    .B(_05055_),
    .Y(_05114_));
 sky130_fd_sc_hd__nand3_2 _11212_ (.A(_05113_),
    .B(_03746_),
    .C(_05114_),
    .Y(_05115_));
 sky130_fd_sc_hd__nand3_1 _11213_ (.A(_05054_),
    .B(_05115_),
    .C(_00820_),
    .Y(_05116_));
 sky130_fd_sc_hd__o21ai_1 _11214_ (.A1(_04830_),
    .A2(_04896_),
    .B1(_05116_),
    .Y(_05117_));
 sky130_fd_sc_hd__nand2_1 _11215_ (.A(_05117_),
    .B(_03281_),
    .Y(_05118_));
 sky130_fd_sc_hd__o211ai_1 _11216_ (.A1(_04830_),
    .A2(_04896_),
    .B1(_03283_),
    .C1(_05116_),
    .Y(_05119_));
 sky130_fd_sc_hd__nand2_1 _11217_ (.A(_05118_),
    .B(_05119_),
    .Y(_05120_));
 sky130_fd_sc_hd__inv_2 _11218_ (.A(_05120_),
    .Y(_05121_));
 sky130_fd_sc_hd__nand3_1 _11219_ (.A(_04824_),
    .B(_04639_),
    .C(_04638_),
    .Y(_05122_));
 sky130_fd_sc_hd__nand2_1 _11220_ (.A(_04820_),
    .B(_04633_),
    .Y(_05123_));
 sky130_fd_sc_hd__inv_2 _11221_ (.A(_04636_),
    .Y(_05124_));
 sky130_fd_sc_hd__nor2_1 _11222_ (.A(_04633_),
    .B(_04820_),
    .Y(_05125_));
 sky130_fd_sc_hd__a21oi_1 _11223_ (.A1(_05123_),
    .A2(_05124_),
    .B1(_05125_),
    .Y(_05126_));
 sky130_fd_sc_hd__nand3_1 _11224_ (.A(_05122_),
    .B(_05126_),
    .C(_04816_),
    .Y(_05127_));
 sky130_fd_sc_hd__nand3_1 _11225_ (.A(_04880_),
    .B(_05121_),
    .C(_05127_),
    .Y(_05128_));
 sky130_fd_sc_hd__nand3_1 _11226_ (.A(_05127_),
    .B(_04878_),
    .C(_03274_),
    .Y(_05129_));
 sky130_fd_sc_hd__nand2_1 _11227_ (.A(_05129_),
    .B(_05120_),
    .Y(_05130_));
 sky130_fd_sc_hd__nand2_1 _11228_ (.A(_05128_),
    .B(_05130_),
    .Y(_05131_));
 sky130_fd_sc_hd__or2_1 _11229_ (.A(_04876_),
    .B(_05131_),
    .X(_05132_));
 sky130_fd_sc_hd__nand2_1 _11230_ (.A(_05131_),
    .B(_04876_),
    .Y(_05133_));
 sky130_fd_sc_hd__clkbuf_4 _11231_ (.A(_00472_),
    .X(_05134_));
 sky130_fd_sc_hd__o21ai_1 _11232_ (.A1(\result_reg_add[12] ),
    .A2(_02649_),
    .B1(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__a31o_1 _11233_ (.A1(_05132_),
    .A2(_02649_),
    .A3(_05133_),
    .B1(_05135_),
    .X(_05136_));
 sky130_fd_sc_hd__inv_2 _11234_ (.A(_05136_),
    .Y(_00256_));
 sky130_fd_sc_hd__nor2_1 _11235_ (.A(_04832_),
    .B(\Oset[2][13] ),
    .Y(_05137_));
 sky130_fd_sc_hd__nor2_1 _11236_ (.A(\Oset[3][13] ),
    .B(_04302_),
    .Y(_05138_));
 sky130_fd_sc_hd__nor2_1 _11237_ (.A(_04832_),
    .B(\Oset[0][13] ),
    .Y(_05139_));
 sky130_fd_sc_hd__o21ai_1 _11238_ (.A1(\Oset[1][13] ),
    .A2(_04302_),
    .B1(_04303_),
    .Y(_05140_));
 sky130_fd_sc_hd__o32a_2 _11239_ (.A1(_04303_),
    .A2(_05137_),
    .A3(_05138_),
    .B1(_05139_),
    .B2(_05140_),
    .X(_05141_));
 sky130_fd_sc_hd__o21ai_1 _11240_ (.A1(_03770_),
    .A2(_05141_),
    .B1(_01156_),
    .Y(_05142_));
 sky130_fd_sc_hd__nor2_1 _11241_ (.A(_04832_),
    .B(\Qset[2][13] ),
    .Y(_05143_));
 sky130_fd_sc_hd__nor2_1 _11242_ (.A(\Qset[3][13] ),
    .B(_04302_),
    .Y(_05144_));
 sky130_fd_sc_hd__nor2_1 _11243_ (.A(_04832_),
    .B(\Qset[0][13] ),
    .Y(_05145_));
 sky130_fd_sc_hd__o21ai_1 _11244_ (.A1(\Qset[1][13] ),
    .A2(_04302_),
    .B1(_04303_),
    .Y(_05146_));
 sky130_fd_sc_hd__o32a_2 _11245_ (.A1(_04303_),
    .A2(_05143_),
    .A3(_05144_),
    .B1(_05145_),
    .B2(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__and2_1 _11246_ (.A(_02458_),
    .B(_02163_),
    .X(_05148_));
 sky130_fd_sc_hd__a211oi_1 _11247_ (.A1(_05147_),
    .A2(_00582_),
    .B1(_03781_),
    .C1(_05148_),
    .Y(_05149_));
 sky130_fd_sc_hd__a2bb2o_1 _11248_ (.A1_N(_05142_),
    .A2_N(_05149_),
    .B1(_00585_),
    .B2(_02466_),
    .X(_05150_));
 sky130_fd_sc_hd__or2_1 _11249_ (.A(_04832_),
    .B(\H[0][13] ),
    .X(_05151_));
 sky130_fd_sc_hd__a21oi_1 _11250_ (.A1(_02469_),
    .A2(_04832_),
    .B1(_04835_),
    .Y(_05152_));
 sky130_fd_sc_hd__mux2_1 _11251_ (.A0(\H[2][13] ),
    .A1(\H[3][13] ),
    .S(_04832_),
    .X(_05153_));
 sky130_fd_sc_hd__a22o_1 _11252_ (.A1(_05151_),
    .A2(_05152_),
    .B1(_05153_),
    .B2(_04835_),
    .X(_05154_));
 sky130_fd_sc_hd__nor2_1 _11253_ (.A(_03758_),
    .B(_05154_),
    .Y(_05155_));
 sky130_fd_sc_hd__a211o_1 _11254_ (.A1(_05150_),
    .A2(_03758_),
    .B1(_00589_),
    .C1(_05155_),
    .X(_05156_));
 sky130_fd_sc_hd__and2_2 _11255_ (.A(_05156_),
    .B(_02473_),
    .X(_05157_));
 sky130_fd_sc_hd__buf_6 _11256_ (.A(_05157_),
    .X(_05158_));
 sky130_fd_sc_hd__a21oi_1 _11257_ (.A1(\Qset[3][13] ),
    .A2(_04857_),
    .B1(_04859_),
    .Y(_05159_));
 sky130_fd_sc_hd__nand2_1 _11258_ (.A(_04855_),
    .B(\Qset[2][13] ),
    .Y(_05160_));
 sky130_fd_sc_hd__a21oi_1 _11259_ (.A1(_04855_),
    .A2(\Qset[0][13] ),
    .B1(_04862_),
    .Y(_05161_));
 sky130_fd_sc_hd__nand2_1 _11260_ (.A(\Qset[1][13] ),
    .B(_04857_),
    .Y(_05162_));
 sky130_fd_sc_hd__a221o_1 _11261_ (.A1(_05159_),
    .A2(_05160_),
    .B1(_05161_),
    .B2(_05162_),
    .C1(_00621_),
    .X(_05163_));
 sky130_fd_sc_hd__a21oi_1 _11262_ (.A1(\Oset[3][13] ),
    .A2(_04857_),
    .B1(_03795_),
    .Y(_05164_));
 sky130_fd_sc_hd__nand2_1 _11263_ (.A(_04415_),
    .B(\Oset[2][13] ),
    .Y(_05165_));
 sky130_fd_sc_hd__a21oi_1 _11264_ (.A1(_04415_),
    .A2(\Oset[0][13] ),
    .B1(_04862_),
    .Y(_05166_));
 sky130_fd_sc_hd__nand2_1 _11265_ (.A(\Oset[1][13] ),
    .B(_04857_),
    .Y(_05167_));
 sky130_fd_sc_hd__a221o_1 _11266_ (.A1(_05164_),
    .A2(_05165_),
    .B1(_05166_),
    .B2(_05167_),
    .C1(_00647_),
    .X(_05168_));
 sky130_fd_sc_hd__a21o_1 _11267_ (.A1(\H[3][13] ),
    .A2(_04857_),
    .B1(_04859_),
    .X(_05169_));
 sky130_fd_sc_hd__a21o_1 _11268_ (.A1(\H[2][13] ),
    .A2(_04855_),
    .B1(_05169_),
    .X(_05170_));
 sky130_fd_sc_hd__a21oi_1 _11269_ (.A1(_04855_),
    .A2(\H[0][13] ),
    .B1(_04862_),
    .Y(_05171_));
 sky130_fd_sc_hd__o21ai_1 _11270_ (.A1(_02469_),
    .A2(_04855_),
    .B1(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__a21oi_1 _11271_ (.A1(_05170_),
    .A2(_05172_),
    .B1(_00626_),
    .Y(_05173_));
 sky130_fd_sc_hd__a311o_2 _11272_ (.A1(_05163_),
    .A2(_05168_),
    .A3(_00626_),
    .B1(_02096_),
    .C1(_05173_),
    .X(_05174_));
 sky130_fd_sc_hd__o21ai_1 _11273_ (.A1(_00820_),
    .A2(_05158_),
    .B1(_05174_),
    .Y(_05175_));
 sky130_fd_sc_hd__nor2_1 _11274_ (.A(_04926_),
    .B(_05158_),
    .Y(_05176_));
 sky130_fd_sc_hd__o21a_1 _11275_ (.A1(_04747_),
    .A2(_04929_),
    .B1(_04932_),
    .X(_05177_));
 sky130_fd_sc_hd__nand2_1 _11276_ (.A(_04690_),
    .B(_04555_),
    .Y(_05178_));
 sky130_fd_sc_hd__nor2_1 _11277_ (.A(_04929_),
    .B(_05178_),
    .Y(_05179_));
 sky130_fd_sc_hd__nand2_1 _11278_ (.A(_05178_),
    .B(_04929_),
    .Y(_05180_));
 sky130_fd_sc_hd__and2b_1 _11279_ (.A_N(_05179_),
    .B(_05180_),
    .X(_05181_));
 sky130_fd_sc_hd__and3_1 _11280_ (.A(_04854_),
    .B(_03079_),
    .C(_03859_),
    .X(_05182_));
 sky130_fd_sc_hd__xnor2_1 _11281_ (.A(_05181_),
    .B(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__nor2_1 _11282_ (.A(_05177_),
    .B(_05183_),
    .Y(_05184_));
 sky130_fd_sc_hd__nand2_1 _11283_ (.A(_05183_),
    .B(_05177_),
    .Y(_05185_));
 sky130_fd_sc_hd__and2b_1 _11284_ (.A_N(_05184_),
    .B(_05185_),
    .X(_05186_));
 sky130_fd_sc_hd__xnor2_1 _11285_ (.A(_05176_),
    .B(_05186_),
    .Y(_05187_));
 sky130_fd_sc_hd__and2_1 _11286_ (.A(_04938_),
    .B(_04935_),
    .X(_05188_));
 sky130_fd_sc_hd__nor2_1 _11287_ (.A(_05187_),
    .B(_05188_),
    .Y(_05189_));
 sky130_fd_sc_hd__inv_2 _11288_ (.A(_05189_),
    .Y(_05190_));
 sky130_fd_sc_hd__nand2_1 _11289_ (.A(_05188_),
    .B(_05187_),
    .Y(_05191_));
 sky130_fd_sc_hd__nand2_1 _11290_ (.A(_05190_),
    .B(_05191_),
    .Y(_05192_));
 sky130_fd_sc_hd__inv_2 _11291_ (.A(_05192_),
    .Y(_05193_));
 sky130_fd_sc_hd__nand2_1 _11292_ (.A(_04944_),
    .B(_04941_),
    .Y(_05194_));
 sky130_fd_sc_hd__or2_1 _11293_ (.A(_05193_),
    .B(_05194_),
    .X(_05195_));
 sky130_fd_sc_hd__nand2_1 _11294_ (.A(_05194_),
    .B(_05193_),
    .Y(_05196_));
 sky130_fd_sc_hd__nand2_1 _11295_ (.A(_05195_),
    .B(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__or2_1 _11296_ (.A(_05026_),
    .B(_05010_),
    .X(_05198_));
 sky130_fd_sc_hd__nand2_1 _11297_ (.A(_05198_),
    .B(_05027_),
    .Y(_05199_));
 sky130_fd_sc_hd__nand2_1 _11298_ (.A(_05197_),
    .B(_05199_),
    .Y(_05200_));
 sky130_fd_sc_hd__nand3b_1 _11299_ (.A_N(_05199_),
    .B(_05195_),
    .C(_05196_),
    .Y(_05201_));
 sky130_fd_sc_hd__nand2_1 _11300_ (.A(_05200_),
    .B(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__inv_2 _11301_ (.A(_05202_),
    .Y(_05203_));
 sky130_fd_sc_hd__nand2_1 _11302_ (.A(_04952_),
    .B(_04947_),
    .Y(_05204_));
 sky130_fd_sc_hd__nand2_1 _11303_ (.A(_05203_),
    .B(_05204_),
    .Y(_05205_));
 sky130_fd_sc_hd__nand3_1 _11304_ (.A(_05202_),
    .B(_04947_),
    .C(_04952_),
    .Y(_05206_));
 sky130_fd_sc_hd__nand2_1 _11305_ (.A(_05205_),
    .B(_05206_),
    .Y(_05207_));
 sky130_fd_sc_hd__a21oi_1 _11306_ (.A1(_04994_),
    .A2(_04997_),
    .B1(_04996_),
    .Y(_05208_));
 sky130_fd_sc_hd__nor2_1 _11307_ (.A(_04973_),
    .B(_04924_),
    .Y(_05209_));
 sky130_fd_sc_hd__nand2_1 _11308_ (.A(_04690_),
    .B(_04982_),
    .Y(_05210_));
 sky130_fd_sc_hd__nor2_1 _11309_ (.A(_04995_),
    .B(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hd__a22o_1 _11310_ (.A1(_04494_),
    .A2(_04982_),
    .B1(_04690_),
    .B2(_04957_),
    .X(_05212_));
 sky130_fd_sc_hd__and2b_1 _11311_ (.A_N(_05211_),
    .B(_05212_),
    .X(_05213_));
 sky130_fd_sc_hd__xnor2_1 _11312_ (.A(_05209_),
    .B(_05213_),
    .Y(_05214_));
 sky130_fd_sc_hd__or2_1 _11313_ (.A(_05208_),
    .B(_05214_),
    .X(_05215_));
 sky130_fd_sc_hd__nand2_1 _11314_ (.A(_05214_),
    .B(_05208_),
    .Y(_05216_));
 sky130_fd_sc_hd__nand2_1 _11315_ (.A(_05215_),
    .B(_05216_),
    .Y(_05217_));
 sky130_fd_sc_hd__or3_1 _11316_ (.A(_04895_),
    .B(_05158_),
    .C(_05217_),
    .X(_05218_));
 sky130_fd_sc_hd__o21ai_1 _11317_ (.A1(_04895_),
    .A2(_05158_),
    .B1(_05217_),
    .Y(_05219_));
 sky130_fd_sc_hd__nand2_1 _11318_ (.A(_05218_),
    .B(_05219_),
    .Y(_05220_));
 sky130_fd_sc_hd__and2b_1 _11319_ (.A_N(_05001_),
    .B(_05004_),
    .X(_05221_));
 sky130_fd_sc_hd__or2_1 _11320_ (.A(_05220_),
    .B(_05221_),
    .X(_05222_));
 sky130_fd_sc_hd__nand2_1 _11321_ (.A(_05221_),
    .B(_05220_),
    .Y(_05223_));
 sky130_fd_sc_hd__nand2_1 _11322_ (.A(_05222_),
    .B(_05223_),
    .Y(_05224_));
 sky130_fd_sc_hd__a21o_1 _11323_ (.A1(_05052_),
    .A2(_05007_),
    .B1(_05224_),
    .X(_05225_));
 sky130_fd_sc_hd__nand3_1 _11324_ (.A(_05052_),
    .B(_05007_),
    .C(_05224_),
    .Y(_05226_));
 sky130_fd_sc_hd__nand3_1 _11325_ (.A(_05225_),
    .B(_03751_),
    .C(_05226_),
    .Y(_05227_));
 sky130_fd_sc_hd__o21ai_1 _11326_ (.A1(_03751_),
    .A2(_05207_),
    .B1(_05227_),
    .Y(_05228_));
 sky130_fd_sc_hd__nand2_1 _11327_ (.A(_05228_),
    .B(_04196_),
    .Y(_05229_));
 sky130_fd_sc_hd__or2_1 _11328_ (.A(_05058_),
    .B(_05110_),
    .X(_05230_));
 sky130_fd_sc_hd__nand2_1 _11329_ (.A(_05114_),
    .B(_05230_),
    .Y(_05231_));
 sky130_fd_sc_hd__nor2_1 _11330_ (.A(_05079_),
    .B(_04309_),
    .Y(_05232_));
 sky130_fd_sc_hd__and2_1 _11331_ (.A(_05070_),
    .B(_05066_),
    .X(_05233_));
 sky130_fd_sc_hd__nor2_1 _11332_ (.A(_03383_),
    .B(_05063_),
    .Y(_05234_));
 sky130_fd_sc_hd__nand2_1 _11333_ (.A(_03652_),
    .B(_03076_),
    .Y(_05235_));
 sky130_fd_sc_hd__nand2_1 _11334_ (.A(_03652_),
    .B(_03110_),
    .Y(_05236_));
 sky130_fd_sc_hd__nand2_1 _11335_ (.A(_05236_),
    .B(_05065_),
    .Y(_05237_));
 sky130_fd_sc_hd__o21a_1 _11336_ (.A1(_05067_),
    .A2(_05235_),
    .B1(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__or2_1 _11337_ (.A(_05234_),
    .B(_05238_),
    .X(_05239_));
 sky130_fd_sc_hd__nand2_1 _11338_ (.A(_05238_),
    .B(_05234_),
    .Y(_05240_));
 sky130_fd_sc_hd__nand2_1 _11339_ (.A(_05239_),
    .B(_05240_),
    .Y(_05241_));
 sky130_fd_sc_hd__nor2_1 _11340_ (.A(_05233_),
    .B(_05241_),
    .Y(_05242_));
 sky130_fd_sc_hd__nand2_1 _11341_ (.A(_05241_),
    .B(_05233_),
    .Y(_05243_));
 sky130_fd_sc_hd__and2b_1 _11342_ (.A_N(_05242_),
    .B(_05243_),
    .X(_05244_));
 sky130_fd_sc_hd__xnor2_1 _11343_ (.A(_05232_),
    .B(_05244_),
    .Y(_05245_));
 sky130_fd_sc_hd__and2_1 _11344_ (.A(_05077_),
    .B(_05074_),
    .X(_05246_));
 sky130_fd_sc_hd__nor2_1 _11345_ (.A(_05245_),
    .B(_05246_),
    .Y(_05247_));
 sky130_fd_sc_hd__inv_2 _11346_ (.A(_05247_),
    .Y(_05248_));
 sky130_fd_sc_hd__nand2_1 _11347_ (.A(_05246_),
    .B(_05245_),
    .Y(_05249_));
 sky130_fd_sc_hd__and2_1 _11348_ (.A(_05248_),
    .B(_05249_),
    .X(_05250_));
 sky130_fd_sc_hd__nand2_1 _11349_ (.A(_05087_),
    .B(_05083_),
    .Y(_05251_));
 sky130_fd_sc_hd__or2_1 _11350_ (.A(_05250_),
    .B(_05251_),
    .X(_05252_));
 sky130_fd_sc_hd__nand2_1 _11351_ (.A(_05251_),
    .B(_05250_),
    .Y(_05253_));
 sky130_fd_sc_hd__nand2_1 _11352_ (.A(_05252_),
    .B(_05253_),
    .Y(_05254_));
 sky130_fd_sc_hd__nor2_1 _11353_ (.A(_05091_),
    .B(_05100_),
    .Y(_05255_));
 sky130_fd_sc_hd__a21oi_1 _11354_ (.A1(_05101_),
    .A2(_05090_),
    .B1(_05255_),
    .Y(_05256_));
 sky130_fd_sc_hd__nor2_1 _11355_ (.A(_04281_),
    .B(_05158_),
    .Y(_05257_));
 sky130_fd_sc_hd__o21a_1 _11356_ (.A1(_05095_),
    .A2(_05094_),
    .B1(_05099_),
    .X(_05258_));
 sky130_fd_sc_hd__nand2_1 _11357_ (.A(_04690_),
    .B(_04651_),
    .Y(_05259_));
 sky130_fd_sc_hd__nand2_1 _11358_ (.A(_04690_),
    .B(_04460_),
    .Y(_05260_));
 sky130_fd_sc_hd__nand2_1 _11359_ (.A(_05260_),
    .B(_05093_),
    .Y(_05261_));
 sky130_fd_sc_hd__o21a_1 _11360_ (.A1(_05094_),
    .A2(_05259_),
    .B1(_05261_),
    .X(_05262_));
 sky130_fd_sc_hd__nor2_1 _11361_ (.A(_04458_),
    .B(_04924_),
    .Y(_05263_));
 sky130_fd_sc_hd__or2_1 _11362_ (.A(_05262_),
    .B(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__nand2_1 _11363_ (.A(_05263_),
    .B(_05262_),
    .Y(_05265_));
 sky130_fd_sc_hd__nand2_1 _11364_ (.A(_05264_),
    .B(_05265_),
    .Y(_05266_));
 sky130_fd_sc_hd__nor2_1 _11365_ (.A(_05258_),
    .B(_05266_),
    .Y(_05267_));
 sky130_fd_sc_hd__nand2_1 _11366_ (.A(_05266_),
    .B(_05258_),
    .Y(_05268_));
 sky130_fd_sc_hd__nor2b_1 _11367_ (.A(_05267_),
    .B_N(_05268_),
    .Y(_05269_));
 sky130_fd_sc_hd__xnor2_1 _11368_ (.A(_05257_),
    .B(_05269_),
    .Y(_05270_));
 sky130_fd_sc_hd__nor2_1 _11369_ (.A(_05256_),
    .B(_05270_),
    .Y(_05271_));
 sky130_fd_sc_hd__inv_2 _11370_ (.A(_05271_),
    .Y(_05272_));
 sky130_fd_sc_hd__nand2_1 _11371_ (.A(_05270_),
    .B(_05256_),
    .Y(_05273_));
 sky130_fd_sc_hd__and2_1 _11372_ (.A(_05272_),
    .B(_05273_),
    .X(_05274_));
 sky130_fd_sc_hd__nand2_1 _11373_ (.A(_05104_),
    .B(_05103_),
    .Y(_05275_));
 sky130_fd_sc_hd__or2_1 _11374_ (.A(_05089_),
    .B(_05102_),
    .X(_05276_));
 sky130_fd_sc_hd__nand2_1 _11375_ (.A(_05275_),
    .B(_05276_),
    .Y(_05277_));
 sky130_fd_sc_hd__or2_1 _11376_ (.A(_05274_),
    .B(_05277_),
    .X(_05278_));
 sky130_fd_sc_hd__nand2_1 _11377_ (.A(_05277_),
    .B(_05274_),
    .Y(_05279_));
 sky130_fd_sc_hd__nand3b_1 _11378_ (.A_N(_05254_),
    .B(_05278_),
    .C(_05279_),
    .Y(_05280_));
 sky130_fd_sc_hd__nand2_1 _11379_ (.A(_05278_),
    .B(_05279_),
    .Y(_05281_));
 sky130_fd_sc_hd__nand2_1 _11380_ (.A(_05281_),
    .B(_05254_),
    .Y(_05282_));
 sky130_fd_sc_hd__nand2_1 _11381_ (.A(_05280_),
    .B(_05282_),
    .Y(_05283_));
 sky130_fd_sc_hd__inv_2 _11382_ (.A(_05283_),
    .Y(_05284_));
 sky130_fd_sc_hd__or2_1 _11383_ (.A(_05088_),
    .B(_05105_),
    .X(_05285_));
 sky130_fd_sc_hd__nand2_1 _11384_ (.A(_05109_),
    .B(_05285_),
    .Y(_05286_));
 sky130_fd_sc_hd__or2_1 _11385_ (.A(_05284_),
    .B(_05286_),
    .X(_05287_));
 sky130_fd_sc_hd__nand2_1 _11386_ (.A(_05286_),
    .B(_05284_),
    .Y(_05288_));
 sky130_fd_sc_hd__nand2_1 _11387_ (.A(_05287_),
    .B(_05288_),
    .Y(_05289_));
 sky130_fd_sc_hd__or2b_1 _11388_ (.A(_04177_),
    .B_N(_04172_),
    .X(_05290_));
 sky130_fd_sc_hd__xor2_1 _11389_ (.A(_04176_),
    .B(_05290_),
    .X(_05291_));
 sky130_fd_sc_hd__nand2_1 _11390_ (.A(_05289_),
    .B(_05291_),
    .Y(_05292_));
 sky130_fd_sc_hd__nand3b_1 _11391_ (.A_N(_05291_),
    .B(_05287_),
    .C(_05288_),
    .Y(_05293_));
 sky130_fd_sc_hd__nand2_1 _11392_ (.A(_05292_),
    .B(_05293_),
    .Y(_05294_));
 sky130_fd_sc_hd__inv_2 _11393_ (.A(_05294_),
    .Y(_05295_));
 sky130_fd_sc_hd__nand2_1 _11394_ (.A(_05231_),
    .B(_05295_),
    .Y(_05296_));
 sky130_fd_sc_hd__nand3_1 _11395_ (.A(_05114_),
    .B(_05294_),
    .C(_05230_),
    .Y(_05297_));
 sky130_fd_sc_hd__nand3_2 _11396_ (.A(_05296_),
    .B(_03746_),
    .C(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hd__nand3_1 _11397_ (.A(_05229_),
    .B(_05298_),
    .C(_00820_),
    .Y(_05299_));
 sky130_fd_sc_hd__o21ai_1 _11398_ (.A1(_00820_),
    .A2(_04974_),
    .B1(_05299_),
    .Y(_05300_));
 sky130_fd_sc_hd__nand2_1 _11399_ (.A(_05300_),
    .B(_02160_),
    .Y(_05301_));
 sky130_fd_sc_hd__o211ai_1 _11400_ (.A1(_04830_),
    .A2(_04974_),
    .B1(_00832_),
    .C1(_05299_),
    .Y(_05302_));
 sky130_fd_sc_hd__nand3b_1 _11401_ (.A_N(_05175_),
    .B(_05301_),
    .C(_05302_),
    .Y(_05303_));
 sky130_fd_sc_hd__nand2_1 _11402_ (.A(_05300_),
    .B(_00832_),
    .Y(_05304_));
 sky130_fd_sc_hd__o211ai_1 _11403_ (.A1(_00820_),
    .A2(_04974_),
    .B1(_02160_),
    .C1(_05299_),
    .Y(_05305_));
 sky130_fd_sc_hd__nand3_1 _11404_ (.A(_05304_),
    .B(_05305_),
    .C(_05175_),
    .Y(_05306_));
 sky130_fd_sc_hd__nand2_1 _11405_ (.A(_05303_),
    .B(_05306_),
    .Y(_05307_));
 sky130_fd_sc_hd__inv_2 _11406_ (.A(_05307_),
    .Y(_05308_));
 sky130_fd_sc_hd__and2_1 _11407_ (.A(_05117_),
    .B(_03296_),
    .X(_05309_));
 sky130_fd_sc_hd__o21bai_1 _11408_ (.A1(_05120_),
    .A2(_05129_),
    .B1_N(_05309_),
    .Y(_05310_));
 sky130_fd_sc_hd__nor2_1 _11409_ (.A(_05308_),
    .B(_05310_),
    .Y(_05311_));
 sky130_fd_sc_hd__inv_2 _11410_ (.A(_05311_),
    .Y(_05312_));
 sky130_fd_sc_hd__nand2_1 _11411_ (.A(_05310_),
    .B(_05308_),
    .Y(_05313_));
 sky130_fd_sc_hd__nand3_2 _11412_ (.A(_05128_),
    .B(_05130_),
    .C(_04876_),
    .Y(_05314_));
 sky130_fd_sc_hd__a21o_1 _11413_ (.A1(_05312_),
    .A2(_05313_),
    .B1(_05314_),
    .X(_05315_));
 sky130_fd_sc_hd__nand3_1 _11414_ (.A(_05312_),
    .B(_05314_),
    .C(_05313_),
    .Y(_05316_));
 sky130_fd_sc_hd__o21ai_1 _11415_ (.A1(\result_reg_add[13] ),
    .A2(_02648_),
    .B1(_05134_),
    .Y(_05317_));
 sky130_fd_sc_hd__a31o_1 _11416_ (.A1(_05315_),
    .A2(_02649_),
    .A3(_05316_),
    .B1(_05317_),
    .X(_05318_));
 sky130_fd_sc_hd__inv_2 _11417_ (.A(_05318_),
    .Y(_00257_));
 sky130_fd_sc_hd__buf_2 _11418_ (.A(_04832_),
    .X(_05319_));
 sky130_fd_sc_hd__nor2_1 _11419_ (.A(_05319_),
    .B(_02483_),
    .Y(_05320_));
 sky130_fd_sc_hd__a211o_1 _11420_ (.A1(_05319_),
    .A2(\Oset[3][14] ),
    .B1(_04303_),
    .C1(_05320_),
    .X(_05321_));
 sky130_fd_sc_hd__nor2_1 _11421_ (.A(_05319_),
    .B(_02486_),
    .Y(_05322_));
 sky130_fd_sc_hd__a211o_1 _11422_ (.A1(_05319_),
    .A2(\Oset[1][14] ),
    .B1(_04835_),
    .C1(_05322_),
    .X(_05323_));
 sky130_fd_sc_hd__nand2_1 _11423_ (.A(_05321_),
    .B(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__nor2_1 _11424_ (.A(_05319_),
    .B(_02476_),
    .Y(_05325_));
 sky130_fd_sc_hd__a211o_1 _11425_ (.A1(_05319_),
    .A2(\Qset[3][14] ),
    .B1(_04303_),
    .C1(_05325_),
    .X(_05326_));
 sky130_fd_sc_hd__nor2_1 _11426_ (.A(_04832_),
    .B(_02479_),
    .Y(_05327_));
 sky130_fd_sc_hd__a211o_1 _11427_ (.A1(_05319_),
    .A2(\Qset[1][14] ),
    .B1(_04835_),
    .C1(_05327_),
    .X(_05328_));
 sky130_fd_sc_hd__nand2_2 _11428_ (.A(_05326_),
    .B(_05328_),
    .Y(_05329_));
 sky130_fd_sc_hd__a21o_1 _11429_ (.A1(_02482_),
    .A2(_02163_),
    .B1(_03781_),
    .X(_05330_));
 sky130_fd_sc_hd__a21o_1 _11430_ (.A1(_00582_),
    .A2(_05329_),
    .B1(_05330_),
    .X(_05331_));
 sky130_fd_sc_hd__o211a_1 _11431_ (.A1(_03770_),
    .A2(_05324_),
    .B1(_01156_),
    .C1(_05331_),
    .X(_05332_));
 sky130_fd_sc_hd__a21o_1 _11432_ (.A1(_00585_),
    .A2(_02489_),
    .B1(_05332_),
    .X(_05333_));
 sky130_fd_sc_hd__or2_1 _11433_ (.A(_05319_),
    .B(\H[0][14] ),
    .X(_05334_));
 sky130_fd_sc_hd__buf_2 _11434_ (.A(_05319_),
    .X(_05335_));
 sky130_fd_sc_hd__a21oi_1 _11435_ (.A1(_02494_),
    .A2(_05335_),
    .B1(_04835_),
    .Y(_05336_));
 sky130_fd_sc_hd__mux2_1 _11436_ (.A0(\H[2][14] ),
    .A1(\H[3][14] ),
    .S(_05319_),
    .X(_05337_));
 sky130_fd_sc_hd__a22o_1 _11437_ (.A1(_05334_),
    .A2(_05336_),
    .B1(_05337_),
    .B2(_04835_),
    .X(_05338_));
 sky130_fd_sc_hd__nor2_1 _11438_ (.A(_03758_),
    .B(_05338_),
    .Y(_05339_));
 sky130_fd_sc_hd__a211o_1 _11439_ (.A1(_05333_),
    .A2(_03758_),
    .B1(_00589_),
    .C1(_05339_),
    .X(_05340_));
 sky130_fd_sc_hd__nand2_4 _11440_ (.A(_05340_),
    .B(_02497_),
    .Y(_05341_));
 sky130_fd_sc_hd__a21o_1 _11441_ (.A1(\H[3][14] ),
    .A2(_04858_),
    .B1(_04859_),
    .X(_05342_));
 sky130_fd_sc_hd__a21o_1 _11442_ (.A1(\H[2][14] ),
    .A2(_04856_),
    .B1(_05342_),
    .X(_05343_));
 sky130_fd_sc_hd__a21oi_1 _11443_ (.A1(_04856_),
    .A2(\H[0][14] ),
    .B1(_04862_),
    .Y(_05344_));
 sky130_fd_sc_hd__o21ai_1 _11444_ (.A1(_02494_),
    .A2(_04856_),
    .B1(_05344_),
    .Y(_05345_));
 sky130_fd_sc_hd__nand2_1 _11445_ (.A(_04855_),
    .B(\Qset[2][14] ),
    .Y(_05346_));
 sky130_fd_sc_hd__a21oi_1 _11446_ (.A1(\Qset[3][14] ),
    .A2(_04857_),
    .B1(_04859_),
    .Y(_05347_));
 sky130_fd_sc_hd__mux2_1 _11447_ (.A0(_02479_),
    .A1(_04053_),
    .S(_03793_),
    .X(_05348_));
 sky130_fd_sc_hd__a221o_1 _11448_ (.A1(_05346_),
    .A2(_05347_),
    .B1(_05348_),
    .B2(_04859_),
    .C1(_00621_),
    .X(_05349_));
 sky130_fd_sc_hd__a21oi_1 _11449_ (.A1(\Oset[3][14] ),
    .A2(_04857_),
    .B1(_04859_),
    .Y(_05350_));
 sky130_fd_sc_hd__nand2_1 _11450_ (.A(_04855_),
    .B(\Oset[2][14] ),
    .Y(_05351_));
 sky130_fd_sc_hd__a21oi_1 _11451_ (.A1(_04855_),
    .A2(\Oset[0][14] ),
    .B1(_04862_),
    .Y(_05352_));
 sky130_fd_sc_hd__nand2_1 _11452_ (.A(\Oset[1][14] ),
    .B(_04858_),
    .Y(_05353_));
 sky130_fd_sc_hd__a221o_1 _11453_ (.A1(_05350_),
    .A2(_05351_),
    .B1(_05352_),
    .B2(_05353_),
    .C1(_00647_),
    .X(_05354_));
 sky130_fd_sc_hd__a21oi_1 _11454_ (.A1(_05349_),
    .A2(_05354_),
    .B1(_01538_),
    .Y(_05355_));
 sky130_fd_sc_hd__a311o_2 _11455_ (.A1(_01538_),
    .A2(_05343_),
    .A3(_05345_),
    .B1(_02096_),
    .C1(_05355_),
    .X(_05356_));
 sky130_fd_sc_hd__o21ai_1 _11456_ (.A1(_04830_),
    .A2(_05341_),
    .B1(_05356_),
    .Y(_05357_));
 sky130_fd_sc_hd__nand2_1 _11457_ (.A(_05296_),
    .B(_05293_),
    .Y(_05358_));
 sky130_fd_sc_hd__nand2_1 _11458_ (.A(_05288_),
    .B(_05280_),
    .Y(_05359_));
 sky130_fd_sc_hd__a21oi_1 _11459_ (.A1(_05243_),
    .A2(_05232_),
    .B1(_05242_),
    .Y(_05360_));
 sky130_fd_sc_hd__nor2_1 _11460_ (.A(_05079_),
    .B(_04495_),
    .Y(_05361_));
 sky130_fd_sc_hd__o21a_1 _11461_ (.A1(_05065_),
    .A2(_05236_),
    .B1(_05240_),
    .X(_05362_));
 sky130_fd_sc_hd__and3_1 _11462_ (.A(_04308_),
    .B(_03745_),
    .C(_03145_),
    .X(_05363_));
 sky130_fd_sc_hd__nand2b_1 _11463_ (.A_N(_05063_),
    .B(_03110_),
    .Y(_05364_));
 sky130_fd_sc_hd__nor2_1 _11464_ (.A(_05235_),
    .B(_05364_),
    .Y(_05365_));
 sky130_fd_sc_hd__nand2_1 _11465_ (.A(_05364_),
    .B(_05235_),
    .Y(_05366_));
 sky130_fd_sc_hd__nor2b_1 _11466_ (.A(_05365_),
    .B_N(_05366_),
    .Y(_05367_));
 sky130_fd_sc_hd__xnor2_1 _11467_ (.A(_05363_),
    .B(_05367_),
    .Y(_05368_));
 sky130_fd_sc_hd__xnor2_1 _11468_ (.A(_05362_),
    .B(_05368_),
    .Y(_05369_));
 sky130_fd_sc_hd__inv_2 _11469_ (.A(_05369_),
    .Y(_05370_));
 sky130_fd_sc_hd__or2_1 _11470_ (.A(_05361_),
    .B(_05370_),
    .X(_05371_));
 sky130_fd_sc_hd__nand2_1 _11471_ (.A(_05370_),
    .B(_05361_),
    .Y(_05372_));
 sky130_fd_sc_hd__nand2_1 _11472_ (.A(_05371_),
    .B(_05372_),
    .Y(_05373_));
 sky130_fd_sc_hd__or2_1 _11473_ (.A(_05360_),
    .B(_05373_),
    .X(_05374_));
 sky130_fd_sc_hd__nand2_1 _11474_ (.A(_05373_),
    .B(_05360_),
    .Y(_05375_));
 sky130_fd_sc_hd__nand2_1 _11475_ (.A(_05374_),
    .B(_05375_),
    .Y(_05376_));
 sky130_fd_sc_hd__nand2_1 _11476_ (.A(_05253_),
    .B(_05248_),
    .Y(_05377_));
 sky130_fd_sc_hd__xor2_1 _11477_ (.A(_05376_),
    .B(_05377_),
    .X(_05378_));
 sky130_fd_sc_hd__inv_2 _11478_ (.A(_05341_),
    .Y(_05379_));
 sky130_fd_sc_hd__nor2_1 _11479_ (.A(_04281_),
    .B(_05379_),
    .Y(_05380_));
 sky130_fd_sc_hd__o21a_1 _11480_ (.A1(_05093_),
    .A2(_05260_),
    .B1(_05265_),
    .X(_05381_));
 sky130_fd_sc_hd__nor2_1 _11481_ (.A(_04458_),
    .B(_05157_),
    .Y(_05382_));
 sky130_fd_sc_hd__nand2_1 _11482_ (.A(_04854_),
    .B(_04460_),
    .Y(_05383_));
 sky130_fd_sc_hd__nor2_1 _11483_ (.A(_05259_),
    .B(_05383_),
    .Y(_05384_));
 sky130_fd_sc_hd__nand2_1 _11484_ (.A(_05383_),
    .B(_05259_),
    .Y(_05385_));
 sky130_fd_sc_hd__nor2b_1 _11485_ (.A(_05384_),
    .B_N(_05385_),
    .Y(_05386_));
 sky130_fd_sc_hd__xnor2_1 _11486_ (.A(_05382_),
    .B(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hd__nor2_1 _11487_ (.A(_05381_),
    .B(_05387_),
    .Y(_05388_));
 sky130_fd_sc_hd__nand2_1 _11488_ (.A(_05387_),
    .B(_05381_),
    .Y(_05389_));
 sky130_fd_sc_hd__nor2b_1 _11489_ (.A(_05388_),
    .B_N(_05389_),
    .Y(_05390_));
 sky130_fd_sc_hd__or2_1 _11490_ (.A(_05380_),
    .B(_05390_),
    .X(_05391_));
 sky130_fd_sc_hd__nand2_1 _11491_ (.A(_05390_),
    .B(_05380_),
    .Y(_05392_));
 sky130_fd_sc_hd__a21o_1 _11492_ (.A1(_05268_),
    .A2(_05257_),
    .B1(_05267_),
    .X(_05393_));
 sky130_fd_sc_hd__a21o_1 _11493_ (.A1(_05391_),
    .A2(_05392_),
    .B1(_05393_),
    .X(_05394_));
 sky130_fd_sc_hd__nand3_1 _11494_ (.A(_05391_),
    .B(_05393_),
    .C(_05392_),
    .Y(_05395_));
 sky130_fd_sc_hd__nand2_1 _11495_ (.A(_05394_),
    .B(_05395_),
    .Y(_05396_));
 sky130_fd_sc_hd__nand2_1 _11496_ (.A(_05279_),
    .B(_05272_),
    .Y(_05397_));
 sky130_fd_sc_hd__xor2_1 _11497_ (.A(_05396_),
    .B(_05397_),
    .X(_05398_));
 sky130_fd_sc_hd__xnor2_1 _11498_ (.A(_05378_),
    .B(_05398_),
    .Y(_05399_));
 sky130_fd_sc_hd__nand2b_1 _11499_ (.A_N(_05359_),
    .B(_05399_),
    .Y(_05400_));
 sky130_fd_sc_hd__a21o_1 _11500_ (.A1(_05288_),
    .A2(_05280_),
    .B1(_05399_),
    .X(_05401_));
 sky130_fd_sc_hd__nand2_1 _11501_ (.A(_05400_),
    .B(_05401_),
    .Y(_05402_));
 sky130_fd_sc_hd__or2b_1 _11502_ (.A(_04163_),
    .B_N(_04180_),
    .X(_05403_));
 sky130_fd_sc_hd__xor2_1 _11503_ (.A(_04178_),
    .B(_05403_),
    .X(_05404_));
 sky130_fd_sc_hd__nand2b_1 _11504_ (.A_N(_05402_),
    .B(_05404_),
    .Y(_05405_));
 sky130_fd_sc_hd__nand2b_1 _11505_ (.A_N(_05404_),
    .B(_05402_),
    .Y(_05406_));
 sky130_fd_sc_hd__nand2_1 _11506_ (.A(_05405_),
    .B(_05406_),
    .Y(_05407_));
 sky130_fd_sc_hd__inv_2 _11507_ (.A(_05407_),
    .Y(_05408_));
 sky130_fd_sc_hd__nand2_1 _11508_ (.A(_05358_),
    .B(_05408_),
    .Y(_05409_));
 sky130_fd_sc_hd__nand3_1 _11509_ (.A(_05407_),
    .B(_05296_),
    .C(_05293_),
    .Y(_05410_));
 sky130_fd_sc_hd__nand3_2 _11510_ (.A(_05409_),
    .B(_05410_),
    .C(_03746_),
    .Y(_05411_));
 sky130_fd_sc_hd__nand2_1 _11511_ (.A(_05225_),
    .B(_05222_),
    .Y(_05412_));
 sky130_fd_sc_hd__nand2_1 _11512_ (.A(_05218_),
    .B(_05215_),
    .Y(_05413_));
 sky130_fd_sc_hd__a21oi_1 _11513_ (.A1(_05209_),
    .A2(_05212_),
    .B1(_05211_),
    .Y(_05414_));
 sky130_fd_sc_hd__nor2_1 _11514_ (.A(_04973_),
    .B(_05158_),
    .Y(_05415_));
 sky130_fd_sc_hd__nand2_1 _11515_ (.A(_04854_),
    .B(_04955_),
    .Y(_05416_));
 sky130_fd_sc_hd__nor2_1 _11516_ (.A(_05210_),
    .B(_05416_),
    .Y(_05417_));
 sky130_fd_sc_hd__nand2_1 _11517_ (.A(_05416_),
    .B(_05210_),
    .Y(_05418_));
 sky130_fd_sc_hd__and2b_1 _11518_ (.A_N(_05417_),
    .B(_05418_),
    .X(_05419_));
 sky130_fd_sc_hd__xnor2_1 _11519_ (.A(_05415_),
    .B(_05419_),
    .Y(_05420_));
 sky130_fd_sc_hd__or2_1 _11520_ (.A(_05414_),
    .B(_05420_),
    .X(_05421_));
 sky130_fd_sc_hd__nand2_1 _11521_ (.A(_05420_),
    .B(_05414_),
    .Y(_05422_));
 sky130_fd_sc_hd__nand2_1 _11522_ (.A(_05421_),
    .B(_05422_),
    .Y(_05423_));
 sky130_fd_sc_hd__or3_1 _11523_ (.A(_04895_),
    .B(_05379_),
    .C(_05423_),
    .X(_05424_));
 sky130_fd_sc_hd__o21ai_1 _11524_ (.A1(_04895_),
    .A2(_05379_),
    .B1(_05423_),
    .Y(_05425_));
 sky130_fd_sc_hd__nand2_1 _11525_ (.A(_05424_),
    .B(_05425_),
    .Y(_05426_));
 sky130_fd_sc_hd__inv_2 _11526_ (.A(_05426_),
    .Y(_05427_));
 sky130_fd_sc_hd__or2_1 _11527_ (.A(_05413_),
    .B(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__nand2_1 _11528_ (.A(_05427_),
    .B(_05413_),
    .Y(_05429_));
 sky130_fd_sc_hd__and2_1 _11529_ (.A(_05428_),
    .B(_05429_),
    .X(_05430_));
 sky130_fd_sc_hd__nand2_1 _11530_ (.A(_05412_),
    .B(_05430_),
    .Y(_05431_));
 sky130_fd_sc_hd__nand3b_1 _11531_ (.A_N(_05430_),
    .B(_05225_),
    .C(_05222_),
    .Y(_05432_));
 sky130_fd_sc_hd__nand3_1 _11532_ (.A(_05431_),
    .B(_05432_),
    .C(_03751_),
    .Y(_05433_));
 sky130_fd_sc_hd__nand2_1 _11533_ (.A(_05205_),
    .B(_05201_),
    .Y(_05434_));
 sky130_fd_sc_hd__nand2_1 _11534_ (.A(_05196_),
    .B(_05190_),
    .Y(_05435_));
 sky130_fd_sc_hd__a21oi_2 _11535_ (.A1(_05185_),
    .A2(_05176_),
    .B1(_05184_),
    .Y(_05436_));
 sky130_fd_sc_hd__nor2_1 _11536_ (.A(_04926_),
    .B(_05379_),
    .Y(_05437_));
 sky130_fd_sc_hd__a21oi_1 _11537_ (.A1(_05182_),
    .A2(_05180_),
    .B1(_05179_),
    .Y(_05438_));
 sky130_fd_sc_hd__nor3_1 _11538_ (.A(_03233_),
    .B(_04345_),
    .C(_05158_),
    .Y(_05439_));
 sky130_fd_sc_hd__nand2_1 _11539_ (.A(_04690_),
    .B(_04744_),
    .Y(_05440_));
 sky130_fd_sc_hd__or3_1 _11540_ (.A(_03051_),
    .B(_04607_),
    .C(_04924_),
    .X(_05441_));
 sky130_fd_sc_hd__nor2_1 _11541_ (.A(_05440_),
    .B(_05441_),
    .Y(_05442_));
 sky130_fd_sc_hd__inv_2 _11542_ (.A(_05442_),
    .Y(_05443_));
 sky130_fd_sc_hd__nand2_1 _11543_ (.A(_05441_),
    .B(_05440_),
    .Y(_05444_));
 sky130_fd_sc_hd__and2_1 _11544_ (.A(_05443_),
    .B(_05444_),
    .X(_05445_));
 sky130_fd_sc_hd__or2_1 _11545_ (.A(_05439_),
    .B(_05445_),
    .X(_05446_));
 sky130_fd_sc_hd__nand2_1 _11546_ (.A(_05445_),
    .B(_05439_),
    .Y(_05447_));
 sky130_fd_sc_hd__nand2_1 _11547_ (.A(_05446_),
    .B(_05447_),
    .Y(_05448_));
 sky130_fd_sc_hd__or2_1 _11548_ (.A(_05438_),
    .B(_05448_),
    .X(_05449_));
 sky130_fd_sc_hd__nand2_1 _11549_ (.A(_05448_),
    .B(_05438_),
    .Y(_05450_));
 sky130_fd_sc_hd__and2_1 _11550_ (.A(_05449_),
    .B(_05450_),
    .X(_05451_));
 sky130_fd_sc_hd__or2_1 _11551_ (.A(_05437_),
    .B(_05451_),
    .X(_05452_));
 sky130_fd_sc_hd__nand2_1 _11552_ (.A(_05451_),
    .B(_05437_),
    .Y(_05453_));
 sky130_fd_sc_hd__nand2_1 _11553_ (.A(_05452_),
    .B(_05453_),
    .Y(_05454_));
 sky130_fd_sc_hd__xnor2_1 _11554_ (.A(_05436_),
    .B(_05454_),
    .Y(_05455_));
 sky130_fd_sc_hd__nand2b_1 _11555_ (.A_N(_05435_),
    .B(_05455_),
    .Y(_05456_));
 sky130_fd_sc_hd__a21o_1 _11556_ (.A1(_05196_),
    .A2(_05190_),
    .B1(_05455_),
    .X(_05457_));
 sky130_fd_sc_hd__nand2_1 _11557_ (.A(_05456_),
    .B(_05457_),
    .Y(_05458_));
 sky130_fd_sc_hd__or2_1 _11558_ (.A(_05041_),
    .B(_05028_),
    .X(_05459_));
 sky130_fd_sc_hd__nand2_1 _11559_ (.A(_05459_),
    .B(_05042_),
    .Y(_05460_));
 sky130_fd_sc_hd__nand2_1 _11560_ (.A(_05458_),
    .B(_05460_),
    .Y(_05461_));
 sky130_fd_sc_hd__nand3b_1 _11561_ (.A_N(_05460_),
    .B(_05456_),
    .C(_05457_),
    .Y(_05462_));
 sky130_fd_sc_hd__nand2_1 _11562_ (.A(_05461_),
    .B(_05462_),
    .Y(_05463_));
 sky130_fd_sc_hd__inv_2 _11563_ (.A(_05463_),
    .Y(_05464_));
 sky130_fd_sc_hd__nand2_1 _11564_ (.A(_05434_),
    .B(_05464_),
    .Y(_05465_));
 sky130_fd_sc_hd__nand3_1 _11565_ (.A(_05463_),
    .B(_05205_),
    .C(_05201_),
    .Y(_05466_));
 sky130_fd_sc_hd__nand3_1 _11566_ (.A(_05465_),
    .B(_05466_),
    .C(_03048_),
    .Y(_05467_));
 sky130_fd_sc_hd__nand2_1 _11567_ (.A(_05433_),
    .B(_05467_),
    .Y(_05468_));
 sky130_fd_sc_hd__nand2_1 _11568_ (.A(_05468_),
    .B(_04196_),
    .Y(_05469_));
 sky130_fd_sc_hd__nand2_1 _11569_ (.A(_05411_),
    .B(_05469_),
    .Y(_05470_));
 sky130_fd_sc_hd__nand2_1 _11570_ (.A(_05470_),
    .B(_04830_),
    .Y(_05471_));
 sky130_fd_sc_hd__nand2_1 _11571_ (.A(_04955_),
    .B(_02096_),
    .Y(_05472_));
 sky130_fd_sc_hd__nand2_1 _11572_ (.A(_05471_),
    .B(_05472_),
    .Y(_05473_));
 sky130_fd_sc_hd__nand2_1 _11573_ (.A(_05473_),
    .B(_02160_),
    .Y(_05474_));
 sky130_fd_sc_hd__nand3_1 _11574_ (.A(_05471_),
    .B(_00832_),
    .C(_05472_),
    .Y(_05475_));
 sky130_fd_sc_hd__nand3b_2 _11575_ (.A_N(_05357_),
    .B(_05474_),
    .C(_05475_),
    .Y(_05476_));
 sky130_fd_sc_hd__nand2_1 _11576_ (.A(_05473_),
    .B(_00832_),
    .Y(_05477_));
 sky130_fd_sc_hd__nand3_1 _11577_ (.A(_05471_),
    .B(_02160_),
    .C(_05472_),
    .Y(_05478_));
 sky130_fd_sc_hd__nand3_1 _11578_ (.A(_05477_),
    .B(_05357_),
    .C(_05478_),
    .Y(_05479_));
 sky130_fd_sc_hd__nand2_1 _11579_ (.A(_05476_),
    .B(_05479_),
    .Y(_05480_));
 sky130_fd_sc_hd__nand2_1 _11580_ (.A(_05480_),
    .B(_05306_),
    .Y(_05481_));
 sky130_fd_sc_hd__nand3b_2 _11581_ (.A_N(_05306_),
    .B(_05476_),
    .C(_05479_),
    .Y(_05482_));
 sky130_fd_sc_hd__nand2_1 _11582_ (.A(_05481_),
    .B(_05482_),
    .Y(_05483_));
 sky130_fd_sc_hd__o21ai_2 _11583_ (.A1(_05314_),
    .A2(_05311_),
    .B1(_05313_),
    .Y(_05484_));
 sky130_fd_sc_hd__or2_1 _11584_ (.A(_05483_),
    .B(_05484_),
    .X(_05485_));
 sky130_fd_sc_hd__nand2_1 _11585_ (.A(_05484_),
    .B(_05483_),
    .Y(_05486_));
 sky130_fd_sc_hd__nand3_1 _11586_ (.A(_05485_),
    .B(_02649_),
    .C(_05486_),
    .Y(_05487_));
 sky130_fd_sc_hd__o21a_1 _11587_ (.A1(\result_reg_add[14] ),
    .A2(_02649_),
    .B1(_01149_),
    .X(_05488_));
 sky130_fd_sc_hd__nand2_1 _11588_ (.A(_05487_),
    .B(_05488_),
    .Y(_05489_));
 sky130_fd_sc_hd__inv_2 _11589_ (.A(_05489_),
    .Y(_00258_));
 sky130_fd_sc_hd__inv_2 _11590_ (.A(_05483_),
    .Y(_05490_));
 sky130_fd_sc_hd__nand2_1 _11591_ (.A(_05484_),
    .B(_05490_),
    .Y(_05491_));
 sky130_fd_sc_hd__nand2_1 _11592_ (.A(_05491_),
    .B(_05482_),
    .Y(_05492_));
 sky130_fd_sc_hd__nand2_1 _11593_ (.A(_05424_),
    .B(_05421_),
    .Y(_05493_));
 sky130_fd_sc_hd__nor2_1 _11594_ (.A(_05335_),
    .B(_02510_),
    .Y(_05494_));
 sky130_fd_sc_hd__nand2_1 _11595_ (.A(_05335_),
    .B(\Oset[1][15] ),
    .Y(_05495_));
 sky130_fd_sc_hd__inv_2 _11596_ (.A(_05495_),
    .Y(_05496_));
 sky130_fd_sc_hd__nor2_1 _11597_ (.A(_05335_),
    .B(_02507_),
    .Y(_05497_));
 sky130_fd_sc_hd__a211o_1 _11598_ (.A1(_05335_),
    .A2(\Oset[3][15] ),
    .B1(_04303_),
    .C1(_05497_),
    .X(_05498_));
 sky130_fd_sc_hd__o31a_1 _11599_ (.A1(_04835_),
    .A2(_05494_),
    .A3(_05496_),
    .B1(_05498_),
    .X(_05499_));
 sky130_fd_sc_hd__inv_2 _11600_ (.A(_05499_),
    .Y(_05500_));
 sky130_fd_sc_hd__a21o_1 _11601_ (.A1(_02506_),
    .A2(_02163_),
    .B1(_03781_),
    .X(_05501_));
 sky130_fd_sc_hd__nand2_1 _11602_ (.A(_04302_),
    .B(_02503_),
    .Y(_05502_));
 sky130_fd_sc_hd__nand2_1 _11603_ (.A(_04076_),
    .B(_05335_),
    .Y(_05503_));
 sky130_fd_sc_hd__o21a_1 _11604_ (.A1(_05335_),
    .A2(\Qset[2][15] ),
    .B1(_04835_),
    .X(_05504_));
 sky130_fd_sc_hd__or2_1 _11605_ (.A(\Qset[3][15] ),
    .B(_04302_),
    .X(_05505_));
 sky130_fd_sc_hd__a32o_1 _11606_ (.A1(_05502_),
    .A2(_05503_),
    .A3(_04303_),
    .B1(_05504_),
    .B2(_05505_),
    .X(_05506_));
 sky130_fd_sc_hd__nor2_1 _11607_ (.A(_02163_),
    .B(_05506_),
    .Y(_05507_));
 sky130_fd_sc_hd__o221a_1 _11608_ (.A1(_03770_),
    .A2(_05500_),
    .B1(_05501_),
    .B2(_05507_),
    .C1(_01156_),
    .X(_05508_));
 sky130_fd_sc_hd__a21oi_1 _11609_ (.A1(_00585_),
    .A2(_02513_),
    .B1(_05508_),
    .Y(_05509_));
 sky130_fd_sc_hd__nor2_1 _11610_ (.A(_05335_),
    .B(_02514_),
    .Y(_05510_));
 sky130_fd_sc_hd__nand2_1 _11611_ (.A(_05335_),
    .B(\H[1][15] ),
    .Y(_05511_));
 sky130_fd_sc_hd__inv_2 _11612_ (.A(_05511_),
    .Y(_05512_));
 sky130_fd_sc_hd__a21o_1 _11613_ (.A1(_05335_),
    .A2(\H[3][15] ),
    .B1(_04303_),
    .X(_05513_));
 sky130_fd_sc_hd__a21o_1 _11614_ (.A1(_04302_),
    .A2(\H[2][15] ),
    .B1(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__o31a_1 _11615_ (.A1(_04835_),
    .A2(_05510_),
    .A3(_05512_),
    .B1(_05514_),
    .X(_05515_));
 sky130_fd_sc_hd__mux2_1 _11616_ (.A0(_05509_),
    .A1(_05515_),
    .S(_03768_),
    .X(_05516_));
 sky130_fd_sc_hd__a21bo_2 _11617_ (.A1(_05516_),
    .A2(_01554_),
    .B1_N(_02519_),
    .X(_05517_));
 sky130_fd_sc_hd__nand2_1 _11618_ (.A(_05517_),
    .B(_04896_),
    .Y(_05518_));
 sky130_fd_sc_hd__a21oi_1 _11619_ (.A1(_05415_),
    .A2(_05418_),
    .B1(_05417_),
    .Y(_05519_));
 sky130_fd_sc_hd__nand2_1 _11620_ (.A(_05341_),
    .B(_04974_),
    .Y(_05520_));
 sky130_fd_sc_hd__nor2_1 _11621_ (.A(_04095_),
    .B(_04924_),
    .Y(_05521_));
 sky130_fd_sc_hd__nor2_1 _11622_ (.A(_04073_),
    .B(_05158_),
    .Y(_05522_));
 sky130_fd_sc_hd__xor2_1 _11623_ (.A(_05521_),
    .B(_05522_),
    .X(_05523_));
 sky130_fd_sc_hd__xor2_1 _11624_ (.A(_05520_),
    .B(_05523_),
    .X(_05524_));
 sky130_fd_sc_hd__xor2_1 _11625_ (.A(_05519_),
    .B(_05524_),
    .X(_05525_));
 sky130_fd_sc_hd__xnor2_1 _11626_ (.A(_05518_),
    .B(_05525_),
    .Y(_05526_));
 sky130_fd_sc_hd__xnor2_1 _11627_ (.A(_05493_),
    .B(_05526_),
    .Y(_05527_));
 sky130_fd_sc_hd__a21oi_1 _11628_ (.A1(_05431_),
    .A2(_05429_),
    .B1(_05527_),
    .Y(_05528_));
 sky130_fd_sc_hd__a31o_1 _11629_ (.A1(_05431_),
    .A2(_05429_),
    .A3(_05527_),
    .B1(_03048_),
    .X(_05529_));
 sky130_fd_sc_hd__nor2_1 _11630_ (.A(_05528_),
    .B(_05529_),
    .Y(_05530_));
 sky130_fd_sc_hd__nor2_1 _11631_ (.A(_03746_),
    .B(_05530_),
    .Y(_05531_));
 sky130_fd_sc_hd__nand2_1 _11632_ (.A(_05465_),
    .B(_05462_),
    .Y(_05532_));
 sky130_fd_sc_hd__o21ai_1 _11633_ (.A1(_05436_),
    .A2(_05454_),
    .B1(_05457_),
    .Y(_05533_));
 sky130_fd_sc_hd__nand2_1 _11634_ (.A(_05341_),
    .B(_03859_),
    .Y(_05534_));
 sky130_fd_sc_hd__or2_1 _11635_ (.A(_03233_),
    .B(_05534_),
    .X(_05535_));
 sky130_fd_sc_hd__nor2_1 _11636_ (.A(_04746_),
    .B(_04924_),
    .Y(_05536_));
 sky130_fd_sc_hd__nor2_1 _11637_ (.A(_04607_),
    .B(_05158_),
    .Y(_05537_));
 sky130_fd_sc_hd__o21a_1 _11638_ (.A1(_05536_),
    .A2(_05537_),
    .B1(_03274_),
    .X(_05538_));
 sky130_fd_sc_hd__nand3_1 _11639_ (.A(_05537_),
    .B(_03274_),
    .C(_05536_),
    .Y(_05539_));
 sky130_fd_sc_hd__nand2_1 _11640_ (.A(_05538_),
    .B(_05539_),
    .Y(_05540_));
 sky130_fd_sc_hd__xnor2_1 _11641_ (.A(_05535_),
    .B(_05540_),
    .Y(_05541_));
 sky130_fd_sc_hd__nand2_1 _11642_ (.A(_05517_),
    .B(_04925_),
    .Y(_05542_));
 sky130_fd_sc_hd__nand2_1 _11643_ (.A(_05447_),
    .B(_05443_),
    .Y(_05543_));
 sky130_fd_sc_hd__xor2_1 _11644_ (.A(_05542_),
    .B(_05543_),
    .X(_05544_));
 sky130_fd_sc_hd__xor2_1 _11645_ (.A(_05541_),
    .B(_05544_),
    .X(_05545_));
 sky130_fd_sc_hd__nand2_1 _11646_ (.A(_05453_),
    .B(_05449_),
    .Y(_05546_));
 sky130_fd_sc_hd__xor2_1 _11647_ (.A(_05545_),
    .B(_05546_),
    .X(_05547_));
 sky130_fd_sc_hd__or2_1 _11648_ (.A(_05047_),
    .B(_05043_),
    .X(_05548_));
 sky130_fd_sc_hd__nand2_1 _11649_ (.A(_05548_),
    .B(_05048_),
    .Y(_05549_));
 sky130_fd_sc_hd__xor2_1 _11650_ (.A(_05547_),
    .B(_05549_),
    .X(_05550_));
 sky130_fd_sc_hd__xor2_1 _11651_ (.A(_05533_),
    .B(_05550_),
    .X(_05551_));
 sky130_fd_sc_hd__xor2_1 _11652_ (.A(_05532_),
    .B(_05551_),
    .X(_05552_));
 sky130_fd_sc_hd__or2_1 _11653_ (.A(_03751_),
    .B(_05552_),
    .X(_05553_));
 sky130_fd_sc_hd__nand2_1 _11654_ (.A(_05531_),
    .B(_05553_),
    .Y(_05554_));
 sky130_fd_sc_hd__nand2_1 _11655_ (.A(_05409_),
    .B(_05405_),
    .Y(_05555_));
 sky130_fd_sc_hd__o21ai_1 _11656_ (.A1(_05378_),
    .A2(_05398_),
    .B1(_05401_),
    .Y(_05556_));
 sky130_fd_sc_hd__or2_1 _11657_ (.A(_04189_),
    .B(_04181_),
    .X(_05557_));
 sky130_fd_sc_hd__and2_1 _11658_ (.A(_05557_),
    .B(_04190_),
    .X(_05558_));
 sky130_fd_sc_hd__o21ai_1 _11659_ (.A1(_05362_),
    .A2(_05368_),
    .B1(_05372_),
    .Y(_05559_));
 sky130_fd_sc_hd__nand2_1 _11660_ (.A(_04690_),
    .B(_05078_),
    .Y(_05560_));
 sky130_fd_sc_hd__a21o_1 _11661_ (.A1(_05366_),
    .A2(_05363_),
    .B1(_05365_),
    .X(_05561_));
 sky130_fd_sc_hd__nand2_1 _11662_ (.A(_04308_),
    .B(_03110_),
    .Y(_05562_));
 sky130_fd_sc_hd__nand2_1 _11663_ (.A(_03790_),
    .B(_03076_),
    .Y(_05563_));
 sky130_fd_sc_hd__xor2_1 _11664_ (.A(_05562_),
    .B(_05563_),
    .X(_05564_));
 sky130_fd_sc_hd__a21oi_1 _11665_ (.A1(_03145_),
    .A2(_04494_),
    .B1(_05564_),
    .Y(_05565_));
 sky130_fd_sc_hd__a31o_1 _11666_ (.A1(_05564_),
    .A2(_03145_),
    .A3(_04494_),
    .B1(_04196_),
    .X(_05566_));
 sky130_fd_sc_hd__nor2_1 _11667_ (.A(_05565_),
    .B(_05566_),
    .Y(_05567_));
 sky130_fd_sc_hd__xor2_1 _11668_ (.A(_05561_),
    .B(_05567_),
    .X(_05568_));
 sky130_fd_sc_hd__xor2_1 _11669_ (.A(_05560_),
    .B(_05568_),
    .X(_05569_));
 sky130_fd_sc_hd__xnor2_1 _11670_ (.A(_05559_),
    .B(_05569_),
    .Y(_05570_));
 sky130_fd_sc_hd__a21bo_1 _11671_ (.A1(_05377_),
    .A2(_05375_),
    .B1_N(_05374_),
    .X(_05571_));
 sky130_fd_sc_hd__xnor2_1 _11672_ (.A(_05570_),
    .B(_05571_),
    .Y(_05572_));
 sky130_fd_sc_hd__a21o_1 _11673_ (.A1(_05389_),
    .A2(_05380_),
    .B1(_05388_),
    .X(_05573_));
 sky130_fd_sc_hd__a21oi_1 _11674_ (.A1(_05382_),
    .A2(_05385_),
    .B1(_05384_),
    .Y(_05574_));
 sky130_fd_sc_hd__nand2_1 _11675_ (.A(_05341_),
    .B(_02734_),
    .Y(_05575_));
 sky130_fd_sc_hd__nand2_1 _11676_ (.A(_05517_),
    .B(_02577_),
    .Y(_05576_));
 sky130_fd_sc_hd__xor2_1 _11677_ (.A(_05575_),
    .B(_05576_),
    .X(_05577_));
 sky130_fd_sc_hd__nand2_1 _11678_ (.A(_04854_),
    .B(_02895_),
    .Y(_05578_));
 sky130_fd_sc_hd__nor2_1 _11679_ (.A(_02897_),
    .B(_05158_),
    .Y(_05579_));
 sky130_fd_sc_hd__xor2_1 _11680_ (.A(_05578_),
    .B(_05579_),
    .X(_05580_));
 sky130_fd_sc_hd__or2_1 _11681_ (.A(_05577_),
    .B(_05580_),
    .X(_05581_));
 sky130_fd_sc_hd__nand2_1 _11682_ (.A(_05580_),
    .B(_05577_),
    .Y(_05582_));
 sky130_fd_sc_hd__a21oi_1 _11683_ (.A1(_05581_),
    .A2(_05582_),
    .B1(_04196_),
    .Y(_05583_));
 sky130_fd_sc_hd__xor2_1 _11684_ (.A(_05574_),
    .B(_05583_),
    .X(_05584_));
 sky130_fd_sc_hd__xor2_1 _11685_ (.A(_05573_),
    .B(_05584_),
    .X(_05585_));
 sky130_fd_sc_hd__a21bo_1 _11686_ (.A1(_05397_),
    .A2(_05394_),
    .B1_N(_05395_),
    .X(_05586_));
 sky130_fd_sc_hd__xor2_1 _11687_ (.A(_05585_),
    .B(_05586_),
    .X(_05587_));
 sky130_fd_sc_hd__xnor2_1 _11688_ (.A(_05572_),
    .B(_05587_),
    .Y(_05588_));
 sky130_fd_sc_hd__xor2_1 _11689_ (.A(_05558_),
    .B(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__xor2_1 _11690_ (.A(_05556_),
    .B(_05589_),
    .X(_05590_));
 sky130_fd_sc_hd__a21oi_1 _11691_ (.A1(_05555_),
    .A2(_05590_),
    .B1(_04196_),
    .Y(_05591_));
 sky130_fd_sc_hd__o21ai_2 _11692_ (.A1(_05555_),
    .A2(_05590_),
    .B1(_05591_),
    .Y(_05592_));
 sky130_fd_sc_hd__nand3_1 _11693_ (.A(_05554_),
    .B(_04830_),
    .C(_05592_),
    .Y(_05593_));
 sky130_fd_sc_hd__nand2_1 _11694_ (.A(_04980_),
    .B(_02096_),
    .Y(_05594_));
 sky130_fd_sc_hd__nand2_1 _11695_ (.A(_05593_),
    .B(_05594_),
    .Y(_05595_));
 sky130_fd_sc_hd__a21o_1 _11696_ (.A1(\H[3][15] ),
    .A2(_04858_),
    .B1(_04859_),
    .X(_05596_));
 sky130_fd_sc_hd__a21o_1 _11697_ (.A1(\H[2][15] ),
    .A2(_04856_),
    .B1(_05596_),
    .X(_05597_));
 sky130_fd_sc_hd__nor2_1 _11698_ (.A(_04858_),
    .B(_02514_),
    .Y(_05598_));
 sky130_fd_sc_hd__a211o_1 _11699_ (.A1(\H[1][15] ),
    .A2(_04858_),
    .B1(_04862_),
    .C1(_05598_),
    .X(_05599_));
 sky130_fd_sc_hd__mux2_1 _11700_ (.A0(\Oset[2][15] ),
    .A1(\Oset[3][15] ),
    .S(_03793_),
    .X(_05600_));
 sky130_fd_sc_hd__nand2_1 _11701_ (.A(\Oset[1][15] ),
    .B(_04857_),
    .Y(_05601_));
 sky130_fd_sc_hd__a21oi_1 _11702_ (.A1(_04415_),
    .A2(\Oset[0][15] ),
    .B1(_03798_),
    .Y(_05602_));
 sky130_fd_sc_hd__a2bb2o_1 _11703_ (.A1_N(_03795_),
    .A2_N(_05600_),
    .B1(_05601_),
    .B2(_05602_),
    .X(_05603_));
 sky130_fd_sc_hd__nand2_1 _11704_ (.A(_04855_),
    .B(\Qset[2][15] ),
    .Y(_05604_));
 sky130_fd_sc_hd__a21oi_1 _11705_ (.A1(\Qset[3][15] ),
    .A2(_04857_),
    .B1(_03795_),
    .Y(_05605_));
 sky130_fd_sc_hd__mux2_1 _11706_ (.A0(_02503_),
    .A1(_04076_),
    .S(_03793_),
    .X(_05606_));
 sky130_fd_sc_hd__a22o_1 _11707_ (.A1(_05604_),
    .A2(_05605_),
    .B1(_05606_),
    .B2(_04859_),
    .X(_05607_));
 sky130_fd_sc_hd__mux2_1 _11708_ (.A0(_05603_),
    .A1(_05607_),
    .S(_00647_),
    .X(_05608_));
 sky130_fd_sc_hd__o21ai_1 _11709_ (.A1(_01538_),
    .A2(_05608_),
    .B1(_00820_),
    .Y(_05609_));
 sky130_fd_sc_hd__a31o_2 _11710_ (.A1(_01538_),
    .A2(_05597_),
    .A3(_05599_),
    .B1(_05609_),
    .X(_05610_));
 sky130_fd_sc_hd__o21ai_1 _11711_ (.A1(_04830_),
    .A2(_05517_),
    .B1(_05610_),
    .Y(_05611_));
 sky130_fd_sc_hd__xor2_1 _11712_ (.A(_00832_),
    .B(_05611_),
    .X(_05612_));
 sky130_fd_sc_hd__nand2_1 _11713_ (.A(_05595_),
    .B(_05612_),
    .Y(_05613_));
 sky130_fd_sc_hd__nand3b_1 _11714_ (.A_N(_05612_),
    .B(_05593_),
    .C(_05594_),
    .Y(_05614_));
 sky130_fd_sc_hd__nand2_1 _11715_ (.A(_05613_),
    .B(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__inv_2 _11716_ (.A(_05476_),
    .Y(_05616_));
 sky130_fd_sc_hd__nand2_1 _11717_ (.A(_05615_),
    .B(_05616_),
    .Y(_05617_));
 sky130_fd_sc_hd__nand3_1 _11718_ (.A(_05613_),
    .B(_05614_),
    .C(_05476_),
    .Y(_05618_));
 sky130_fd_sc_hd__nand2_1 _11719_ (.A(_05617_),
    .B(_05618_),
    .Y(_05619_));
 sky130_fd_sc_hd__inv_2 _11720_ (.A(_05619_),
    .Y(_05620_));
 sky130_fd_sc_hd__nand2_1 _11721_ (.A(_05492_),
    .B(_05620_),
    .Y(_05621_));
 sky130_fd_sc_hd__nand3_1 _11722_ (.A(_05491_),
    .B(_05482_),
    .C(_05619_),
    .Y(_05622_));
 sky130_fd_sc_hd__nand3_1 _11723_ (.A(_05621_),
    .B(_02649_),
    .C(_05622_),
    .Y(_05623_));
 sky130_fd_sc_hd__o21a_1 _11724_ (.A1(\result_reg_add[15] ),
    .A2(_02649_),
    .B1(_01149_),
    .X(_05624_));
 sky130_fd_sc_hd__nand2_1 _11725_ (.A(_05623_),
    .B(_05624_),
    .Y(_05625_));
 sky130_fd_sc_hd__inv_2 _11726_ (.A(_05625_),
    .Y(_00259_));
 sky130_fd_sc_hd__or3_1 _11727_ (.A(CMD_addition),
    .B(_00832_),
    .C(_06269_),
    .X(_05626_));
 sky130_fd_sc_hd__clkbuf_4 _11728_ (.A(_05626_),
    .X(_05627_));
 sky130_fd_sc_hd__buf_6 _11729_ (.A(_05627_),
    .X(_05628_));
 sky130_fd_sc_hd__a21oi_1 _11730_ (.A1(_05628_),
    .A2(_00610_),
    .B1(_02650_),
    .Y(_05629_));
 sky130_fd_sc_hd__o21ai_1 _11731_ (.A1(_05628_),
    .A2(_02645_),
    .B1(_05629_),
    .Y(_05630_));
 sky130_fd_sc_hd__inv_2 _11732_ (.A(_05630_),
    .Y(_00260_));
 sky130_fd_sc_hd__clkbuf_4 _11733_ (.A(_05627_),
    .X(_05631_));
 sky130_fd_sc_hd__nor2_1 _11734_ (.A(_05631_),
    .B(_02750_),
    .Y(_05632_));
 sky130_fd_sc_hd__a211o_1 _11735_ (.A1(_00702_),
    .A2(_05628_),
    .B1(_02753_),
    .C1(_05632_),
    .X(_05633_));
 sky130_fd_sc_hd__inv_2 _11736_ (.A(_05633_),
    .Y(_00261_));
 sky130_fd_sc_hd__clkbuf_4 _11737_ (.A(_00635_),
    .X(_05634_));
 sky130_fd_sc_hd__nor2_1 _11738_ (.A(_05631_),
    .B(_02860_),
    .Y(_05635_));
 sky130_fd_sc_hd__a211o_1 _11739_ (.A1(_00728_),
    .A2(_05628_),
    .B1(_05634_),
    .C1(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__inv_2 _11740_ (.A(_05636_),
    .Y(_00262_));
 sky130_fd_sc_hd__nor2_1 _11741_ (.A(_05631_),
    .B(_02986_),
    .Y(_05637_));
 sky130_fd_sc_hd__a211o_1 _11742_ (.A1(_00770_),
    .A2(_05631_),
    .B1(_05634_),
    .C1(_05637_),
    .X(_05638_));
 sky130_fd_sc_hd__inv_2 _11743_ (.A(_05638_),
    .Y(_00263_));
 sky130_fd_sc_hd__nor2_1 _11744_ (.A(_05627_),
    .B(_03293_),
    .Y(_05639_));
 sky130_fd_sc_hd__a211o_1 _11745_ (.A1(_00788_),
    .A2(_05631_),
    .B1(_05634_),
    .C1(_05639_),
    .X(_05640_));
 sky130_fd_sc_hd__inv_2 _11746_ (.A(_05640_),
    .Y(_00264_));
 sky130_fd_sc_hd__nor2_1 _11747_ (.A(_05627_),
    .B(_03449_),
    .Y(_05641_));
 sky130_fd_sc_hd__a211o_1 _11748_ (.A1(_00841_),
    .A2(_05631_),
    .B1(_05634_),
    .C1(_05641_),
    .X(_05642_));
 sky130_fd_sc_hd__inv_2 _11749_ (.A(_05642_),
    .Y(_00265_));
 sky130_fd_sc_hd__nor2_1 _11750_ (.A(_05627_),
    .B(_03601_),
    .Y(_05643_));
 sky130_fd_sc_hd__a211o_1 _11751_ (.A1(_00865_),
    .A2(_05631_),
    .B1(_05634_),
    .C1(_05643_),
    .X(_05644_));
 sky130_fd_sc_hd__inv_2 _11752_ (.A(_05644_),
    .Y(_00266_));
 sky130_fd_sc_hd__nor2_1 _11753_ (.A(_05627_),
    .B(_03740_),
    .Y(_05645_));
 sky130_fd_sc_hd__a211o_1 _11754_ (.A1(_00883_),
    .A2(_05631_),
    .B1(_05634_),
    .C1(_05645_),
    .X(_05646_));
 sky130_fd_sc_hd__inv_2 _11755_ (.A(_05646_),
    .Y(_00267_));
 sky130_fd_sc_hd__a21oi_1 _11756_ (.A1(_05628_),
    .A2(_00912_),
    .B1(_02650_),
    .Y(_05647_));
 sky130_fd_sc_hd__o21ai_1 _11757_ (.A1(_05628_),
    .A2(_04256_),
    .B1(_05647_),
    .Y(_05648_));
 sky130_fd_sc_hd__inv_2 _11758_ (.A(_05648_),
    .Y(_00268_));
 sky130_fd_sc_hd__nor2_1 _11759_ (.A(_05627_),
    .B(_04444_),
    .Y(_05649_));
 sky130_fd_sc_hd__a211o_1 _11760_ (.A1(_00932_),
    .A2(_05631_),
    .B1(_05634_),
    .C1(_05649_),
    .X(_05650_));
 sky130_fd_sc_hd__inv_2 _11761_ (.A(_05650_),
    .Y(_00269_));
 sky130_fd_sc_hd__nor2_1 _11762_ (.A(_05627_),
    .B(_04642_),
    .Y(_05651_));
 sky130_fd_sc_hd__a211o_1 _11763_ (.A1(_00958_),
    .A2(_05631_),
    .B1(_05634_),
    .C1(_05651_),
    .X(_05652_));
 sky130_fd_sc_hd__inv_2 _11764_ (.A(_05652_),
    .Y(_00270_));
 sky130_fd_sc_hd__a21oi_1 _11765_ (.A1(_05628_),
    .A2(_00991_),
    .B1(_02650_),
    .Y(_05653_));
 sky130_fd_sc_hd__o21ai_1 _11766_ (.A1(_05628_),
    .A2(_04826_),
    .B1(_05653_),
    .Y(_05654_));
 sky130_fd_sc_hd__inv_2 _11767_ (.A(_05654_),
    .Y(_00271_));
 sky130_fd_sc_hd__inv_2 _11768_ (.A(_05626_),
    .Y(_05655_));
 sky130_fd_sc_hd__a21o_1 _11769_ (.A1(_05627_),
    .A2(_01016_),
    .B1(_02115_),
    .X(_05656_));
 sky130_fd_sc_hd__a31o_1 _11770_ (.A1(_05132_),
    .A2(_05133_),
    .A3(_05655_),
    .B1(_05656_),
    .X(_05657_));
 sky130_fd_sc_hd__inv_2 _11771_ (.A(_05657_),
    .Y(_00272_));
 sky130_fd_sc_hd__a21o_1 _11772_ (.A1(_05627_),
    .A2(_01035_),
    .B1(_02115_),
    .X(_05658_));
 sky130_fd_sc_hd__a31o_1 _11773_ (.A1(_05315_),
    .A2(_05316_),
    .A3(_05655_),
    .B1(_05658_),
    .X(_05659_));
 sky130_fd_sc_hd__inv_2 _11774_ (.A(_05659_),
    .Y(_00273_));
 sky130_fd_sc_hd__nand3_1 _11775_ (.A(_05485_),
    .B(_05486_),
    .C(_05655_),
    .Y(_05660_));
 sky130_fd_sc_hd__a21oi_1 _11776_ (.A1(_05628_),
    .A2(_01067_),
    .B1(_02650_),
    .Y(_05661_));
 sky130_fd_sc_hd__nand2_1 _11777_ (.A(_05660_),
    .B(_05661_),
    .Y(_05662_));
 sky130_fd_sc_hd__inv_2 _11778_ (.A(_05662_),
    .Y(_00274_));
 sky130_fd_sc_hd__nand3_1 _11779_ (.A(_05621_),
    .B(_05622_),
    .C(_05655_),
    .Y(_05663_));
 sky130_fd_sc_hd__a21oi_1 _11780_ (.A1(_05628_),
    .A2(_01093_),
    .B1(_02650_),
    .Y(_05664_));
 sky130_fd_sc_hd__nand2_1 _11781_ (.A(_05663_),
    .B(_05664_),
    .Y(_05665_));
 sky130_fd_sc_hd__inv_2 _11782_ (.A(_05665_),
    .Y(_00275_));
 sky130_fd_sc_hd__inv_2 _11783_ (.A(_02093_),
    .Y(_05666_));
 sky130_fd_sc_hd__nor2_2 _11784_ (.A(_06269_),
    .B(_05666_),
    .Y(_05667_));
 sky130_fd_sc_hd__inv_2 _11785_ (.A(_05667_),
    .Y(_05668_));
 sky130_fd_sc_hd__nor2_4 _11786_ (.A(_00528_),
    .B(_05668_),
    .Y(_05669_));
 sky130_fd_sc_hd__clkbuf_4 _11787_ (.A(_05669_),
    .X(_05670_));
 sky130_fd_sc_hd__nand2_1 _11788_ (.A(_02621_),
    .B(_05670_),
    .Y(_05671_));
 sky130_fd_sc_hd__o211a_1 _11789_ (.A1(\result_reg_mul[0] ),
    .A2(_05670_),
    .B1(_02105_),
    .C1(_05671_),
    .X(_00276_));
 sky130_fd_sc_hd__buf_4 _11790_ (.A(_01148_),
    .X(_05672_));
 sky130_fd_sc_hd__inv_2 _11791_ (.A(_05669_),
    .Y(_05673_));
 sky130_fd_sc_hd__a21o_1 _11792_ (.A1(_02737_),
    .A2(_02740_),
    .B1(_05673_),
    .X(_05674_));
 sky130_fd_sc_hd__o211a_1 _11793_ (.A1(\result_reg_mul[1] ),
    .A2(_05670_),
    .B1(_05672_),
    .C1(_05674_),
    .X(_00277_));
 sky130_fd_sc_hd__a21o_1 _11794_ (.A1(_02828_),
    .A2(_02830_),
    .B1(_05673_),
    .X(_05675_));
 sky130_fd_sc_hd__o211a_1 _11795_ (.A1(\result_reg_mul[2] ),
    .A2(_05670_),
    .B1(_05672_),
    .C1(_05675_),
    .X(_00278_));
 sky130_fd_sc_hd__nand2_1 _11796_ (.A(_02957_),
    .B(_05670_),
    .Y(_05676_));
 sky130_fd_sc_hd__o211a_1 _11797_ (.A1(\result_reg_mul[3] ),
    .A2(_05670_),
    .B1(_05672_),
    .C1(_05676_),
    .X(_00279_));
 sky130_fd_sc_hd__clkbuf_4 _11798_ (.A(_05669_),
    .X(_05677_));
 sky130_fd_sc_hd__o21ai_1 _11799_ (.A1(\result_reg_mul[4] ),
    .A2(_05677_),
    .B1(_05134_),
    .Y(_05678_));
 sky130_fd_sc_hd__a31o_1 _11800_ (.A1(_03234_),
    .A2(_03276_),
    .A3(_05670_),
    .B1(_05678_),
    .X(_05679_));
 sky130_fd_sc_hd__inv_2 _11801_ (.A(_05679_),
    .Y(_00280_));
 sky130_fd_sc_hd__o21ai_1 _11802_ (.A1(\result_reg_mul[5] ),
    .A2(_05677_),
    .B1(_05134_),
    .Y(_05680_));
 sky130_fd_sc_hd__a31o_1 _11803_ (.A1(_03416_),
    .A2(_03417_),
    .A3(_05670_),
    .B1(_05680_),
    .X(_05681_));
 sky130_fd_sc_hd__inv_2 _11804_ (.A(_05681_),
    .Y(_00281_));
 sky130_fd_sc_hd__clkbuf_4 _11805_ (.A(_00472_),
    .X(_05682_));
 sky130_fd_sc_hd__o21ai_1 _11806_ (.A1(\result_reg_mul[6] ),
    .A2(_05669_),
    .B1(_05682_),
    .Y(_05683_));
 sky130_fd_sc_hd__a31o_1 _11807_ (.A1(_03569_),
    .A2(_03570_),
    .A3(_05677_),
    .B1(_05683_),
    .X(_05684_));
 sky130_fd_sc_hd__inv_2 _11808_ (.A(_05684_),
    .Y(_00282_));
 sky130_fd_sc_hd__o21ai_1 _11809_ (.A1(\result_reg_mul[7] ),
    .A2(_05669_),
    .B1(_05682_),
    .Y(_05685_));
 sky130_fd_sc_hd__a31o_1 _11810_ (.A1(_03682_),
    .A2(_03704_),
    .A3(_05677_),
    .B1(_05685_),
    .X(_05686_));
 sky130_fd_sc_hd__inv_2 _11811_ (.A(_05686_),
    .Y(_00283_));
 sky130_fd_sc_hd__o21ai_1 _11812_ (.A1(\result_reg_mul[8] ),
    .A2(_05669_),
    .B1(_05682_),
    .Y(_05687_));
 sky130_fd_sc_hd__a31o_1 _11813_ (.A1(_04198_),
    .A2(_04248_),
    .A3(_05677_),
    .B1(_05687_),
    .X(_05688_));
 sky130_fd_sc_hd__inv_2 _11814_ (.A(_05688_),
    .Y(_00284_));
 sky130_fd_sc_hd__o21ai_1 _11815_ (.A1(\result_reg_mul[9] ),
    .A2(_05669_),
    .B1(_05682_),
    .Y(_05689_));
 sky130_fd_sc_hd__a31o_1 _11816_ (.A1(_04408_),
    .A2(_04409_),
    .A3(_05677_),
    .B1(_05689_),
    .X(_05690_));
 sky130_fd_sc_hd__inv_2 _11817_ (.A(_05690_),
    .Y(_00285_));
 sky130_fd_sc_hd__o21ai_1 _11818_ (.A1(\result_reg_mul[10] ),
    .A2(_05669_),
    .B1(_05682_),
    .Y(_05691_));
 sky130_fd_sc_hd__a31o_1 _11819_ (.A1(_04527_),
    .A2(_04605_),
    .A3(_05677_),
    .B1(_05691_),
    .X(_05692_));
 sky130_fd_sc_hd__inv_2 _11820_ (.A(_05692_),
    .Y(_00286_));
 sky130_fd_sc_hd__a21o_1 _11821_ (.A1(_04722_),
    .A2(_04791_),
    .B1(_05673_),
    .X(_05693_));
 sky130_fd_sc_hd__o211a_1 _11822_ (.A1(\result_reg_mul[11] ),
    .A2(_05670_),
    .B1(_05672_),
    .C1(_05693_),
    .X(_00287_));
 sky130_fd_sc_hd__o21ai_1 _11823_ (.A1(\result_reg_mul[12] ),
    .A2(_05669_),
    .B1(_05682_),
    .Y(_05694_));
 sky130_fd_sc_hd__a31o_1 _11824_ (.A1(_05054_),
    .A2(_05115_),
    .A3(_05677_),
    .B1(_05694_),
    .X(_05695_));
 sky130_fd_sc_hd__inv_2 _11825_ (.A(_05695_),
    .Y(_00288_));
 sky130_fd_sc_hd__o21ai_1 _11826_ (.A1(\result_reg_mul[13] ),
    .A2(_05669_),
    .B1(_05682_),
    .Y(_05696_));
 sky130_fd_sc_hd__a31o_1 _11827_ (.A1(_05229_),
    .A2(_05298_),
    .A3(_05677_),
    .B1(_05696_),
    .X(_05697_));
 sky130_fd_sc_hd__inv_2 _11828_ (.A(_05697_),
    .Y(_00289_));
 sky130_fd_sc_hd__o21a_1 _11829_ (.A1(\result_reg_mul[14] ),
    .A2(_05677_),
    .B1(_01149_),
    .X(_05698_));
 sky130_fd_sc_hd__o21ai_1 _11830_ (.A1(_05673_),
    .A2(_05470_),
    .B1(_05698_),
    .Y(_05699_));
 sky130_fd_sc_hd__inv_2 _11831_ (.A(_05699_),
    .Y(_00290_));
 sky130_fd_sc_hd__a21o_1 _11832_ (.A1(_05554_),
    .A2(_05592_),
    .B1(_05673_),
    .X(_05700_));
 sky130_fd_sc_hd__o211a_1 _11833_ (.A1(\result_reg_mul[15] ),
    .A2(_05670_),
    .B1(_05672_),
    .C1(_05700_),
    .X(_00291_));
 sky130_fd_sc_hd__and3_1 _11834_ (.A(_05667_),
    .B(_04830_),
    .C(_00528_),
    .X(_05701_));
 sky130_fd_sc_hd__buf_4 _11835_ (.A(_05701_),
    .X(_05702_));
 sky130_fd_sc_hd__buf_4 _11836_ (.A(_05702_),
    .X(_05703_));
 sky130_fd_sc_hd__nor2_1 _11837_ (.A(\result_reg_mac[0] ),
    .B(_05702_),
    .Y(_05704_));
 sky130_fd_sc_hd__a211o_1 _11838_ (.A1(_02646_),
    .A2(_05703_),
    .B1(_05634_),
    .C1(_05704_),
    .X(_05705_));
 sky130_fd_sc_hd__inv_2 _11839_ (.A(_05705_),
    .Y(_00292_));
 sky130_fd_sc_hd__inv_2 _11840_ (.A(_05702_),
    .Y(_05706_));
 sky130_fd_sc_hd__buf_4 _11841_ (.A(_05706_),
    .X(_05707_));
 sky130_fd_sc_hd__nor2_1 _11842_ (.A(_05706_),
    .B(_02750_),
    .Y(_05708_));
 sky130_fd_sc_hd__a211o_1 _11843_ (.A1(_00694_),
    .A2(_05707_),
    .B1(_05634_),
    .C1(_05708_),
    .X(_05709_));
 sky130_fd_sc_hd__inv_2 _11844_ (.A(_05709_),
    .Y(_00293_));
 sky130_fd_sc_hd__buf_4 _11845_ (.A(_00635_),
    .X(_05710_));
 sky130_fd_sc_hd__nor2_1 _11846_ (.A(_05706_),
    .B(_02860_),
    .Y(_05711_));
 sky130_fd_sc_hd__a211o_1 _11847_ (.A1(_00724_),
    .A2(_05707_),
    .B1(_05710_),
    .C1(_05711_),
    .X(_05712_));
 sky130_fd_sc_hd__inv_2 _11848_ (.A(_05712_),
    .Y(_00294_));
 sky130_fd_sc_hd__nor2_1 _11849_ (.A(_05706_),
    .B(_02986_),
    .Y(_05713_));
 sky130_fd_sc_hd__a211o_1 _11850_ (.A1(_00761_),
    .A2(_05707_),
    .B1(_05710_),
    .C1(_05713_),
    .X(_05714_));
 sky130_fd_sc_hd__inv_2 _11851_ (.A(_05714_),
    .Y(_00295_));
 sky130_fd_sc_hd__nor2_1 _11852_ (.A(_05706_),
    .B(_03293_),
    .Y(_05715_));
 sky130_fd_sc_hd__a211o_1 _11853_ (.A1(_00785_),
    .A2(_05707_),
    .B1(_05710_),
    .C1(_05715_),
    .X(_05716_));
 sky130_fd_sc_hd__inv_2 _11854_ (.A(_05716_),
    .Y(_00296_));
 sky130_fd_sc_hd__nor2_1 _11855_ (.A(_05706_),
    .B(_03449_),
    .Y(_05717_));
 sky130_fd_sc_hd__a211o_1 _11856_ (.A1(_00811_),
    .A2(_05707_),
    .B1(_05710_),
    .C1(_05717_),
    .X(_05718_));
 sky130_fd_sc_hd__inv_2 _11857_ (.A(_05718_),
    .Y(_00297_));
 sky130_fd_sc_hd__nor2_1 _11858_ (.A(_05706_),
    .B(_03601_),
    .Y(_05719_));
 sky130_fd_sc_hd__a211o_1 _11859_ (.A1(_00856_),
    .A2(_05707_),
    .B1(_05710_),
    .C1(_05719_),
    .X(_05720_));
 sky130_fd_sc_hd__inv_2 _11860_ (.A(_05720_),
    .Y(_00298_));
 sky130_fd_sc_hd__nor2_1 _11861_ (.A(_05706_),
    .B(_03740_),
    .Y(_05721_));
 sky130_fd_sc_hd__a211o_1 _11862_ (.A1(_00880_),
    .A2(_05707_),
    .B1(_05710_),
    .C1(_05721_),
    .X(_05722_));
 sky130_fd_sc_hd__inv_2 _11863_ (.A(_05722_),
    .Y(_00299_));
 sky130_fd_sc_hd__nor2_1 _11864_ (.A(\result_reg_mac[8] ),
    .B(_05702_),
    .Y(_05723_));
 sky130_fd_sc_hd__a211o_1 _11865_ (.A1(_04257_),
    .A2(_05703_),
    .B1(_05710_),
    .C1(_05723_),
    .X(_05724_));
 sky130_fd_sc_hd__inv_2 _11866_ (.A(_05724_),
    .Y(_00300_));
 sky130_fd_sc_hd__nor2_1 _11867_ (.A(_05706_),
    .B(_04444_),
    .Y(_05725_));
 sky130_fd_sc_hd__a211o_1 _11868_ (.A1(_00929_),
    .A2(_05707_),
    .B1(_05710_),
    .C1(_05725_),
    .X(_05726_));
 sky130_fd_sc_hd__inv_2 _11869_ (.A(_05726_),
    .Y(_00301_));
 sky130_fd_sc_hd__nor2_1 _11870_ (.A(_05706_),
    .B(_04642_),
    .Y(_05727_));
 sky130_fd_sc_hd__a211o_1 _11871_ (.A1(_00955_),
    .A2(_05707_),
    .B1(_05710_),
    .C1(_05727_),
    .X(_05728_));
 sky130_fd_sc_hd__inv_2 _11872_ (.A(_05728_),
    .Y(_00302_));
 sky130_fd_sc_hd__o21a_1 _11873_ (.A1(\result_reg_mac[11] ),
    .A2(_05703_),
    .B1(_01149_),
    .X(_05729_));
 sky130_fd_sc_hd__o21ai_1 _11874_ (.A1(_05707_),
    .A2(_04826_),
    .B1(_05729_),
    .Y(_05730_));
 sky130_fd_sc_hd__inv_2 _11875_ (.A(_05730_),
    .Y(_00303_));
 sky130_fd_sc_hd__o21ai_1 _11876_ (.A1(\result_reg_mac[12] ),
    .A2(_05703_),
    .B1(_05682_),
    .Y(_05731_));
 sky130_fd_sc_hd__a31o_1 _11877_ (.A1(_05132_),
    .A2(_05133_),
    .A3(_05703_),
    .B1(_05731_),
    .X(_05732_));
 sky130_fd_sc_hd__inv_2 _11878_ (.A(_05732_),
    .Y(_00304_));
 sky130_fd_sc_hd__o21ai_1 _11879_ (.A1(\result_reg_mac[13] ),
    .A2(_05702_),
    .B1(_05682_),
    .Y(_05733_));
 sky130_fd_sc_hd__a31o_1 _11880_ (.A1(_05315_),
    .A2(_05316_),
    .A3(_05703_),
    .B1(_05733_),
    .X(_05734_));
 sky130_fd_sc_hd__inv_2 _11881_ (.A(_05734_),
    .Y(_00305_));
 sky130_fd_sc_hd__nand3_1 _11882_ (.A(_05485_),
    .B(_05486_),
    .C(_05703_),
    .Y(_05735_));
 sky130_fd_sc_hd__o21a_1 _11883_ (.A1(\result_reg_mac[14] ),
    .A2(_05703_),
    .B1(_01149_),
    .X(_05736_));
 sky130_fd_sc_hd__nand2_1 _11884_ (.A(_05735_),
    .B(_05736_),
    .Y(_05737_));
 sky130_fd_sc_hd__inv_2 _11885_ (.A(_05737_),
    .Y(_00306_));
 sky130_fd_sc_hd__nand3_1 _11886_ (.A(_05621_),
    .B(_05622_),
    .C(_05703_),
    .Y(_05738_));
 sky130_fd_sc_hd__o21a_1 _11887_ (.A1(\result_reg_mac[15] ),
    .A2(_05703_),
    .B1(_01149_),
    .X(_05739_));
 sky130_fd_sc_hd__nand2_1 _11888_ (.A(_05738_),
    .B(_05739_),
    .Y(_05740_));
 sky130_fd_sc_hd__inv_2 _11889_ (.A(_05740_),
    .Y(_00307_));
 sky130_fd_sc_hd__nor2_2 _11890_ (.A(_05668_),
    .B(_01602_),
    .Y(_05741_));
 sky130_fd_sc_hd__or3_1 _11891_ (.A(_00659_),
    .B(_02115_),
    .C(_05741_),
    .X(_05742_));
 sky130_fd_sc_hd__inv_2 _11892_ (.A(_05742_),
    .Y(_00308_));
 sky130_fd_sc_hd__clkbuf_4 _11893_ (.A(_05741_),
    .X(_05743_));
 sky130_fd_sc_hd__clkbuf_4 _11894_ (.A(_00590_),
    .X(_05744_));
 sky130_fd_sc_hd__clkbuf_4 _11895_ (.A(_01158_),
    .X(_05745_));
 sky130_fd_sc_hd__inv_2 _11896_ (.A(_02570_),
    .Y(_05746_));
 sky130_fd_sc_hd__nor2_1 _11897_ (.A(_01554_),
    .B(_05746_),
    .Y(_05747_));
 sky130_fd_sc_hd__a221o_2 _11898_ (.A1(_05744_),
    .A2(_02538_),
    .B1(_05745_),
    .B2(_02550_),
    .C1(_05747_),
    .X(_05748_));
 sky130_fd_sc_hd__clkbuf_4 _11899_ (.A(_00589_),
    .X(_05749_));
 sky130_fd_sc_hd__nand2_2 _11900_ (.A(_02790_),
    .B(_02793_),
    .Y(_05750_));
 sky130_fd_sc_hd__inv_2 _11901_ (.A(_05750_),
    .Y(_05751_));
 sky130_fd_sc_hd__nor2_1 _11902_ (.A(_00591_),
    .B(_05751_),
    .Y(_05752_));
 sky130_fd_sc_hd__a221o_2 _11903_ (.A1(_01158_),
    .A2(_02807_),
    .B1(_02817_),
    .B2(_05749_),
    .C1(_05752_),
    .X(_05753_));
 sky130_fd_sc_hd__inv_2 _11904_ (.A(_02118_),
    .Y(_05754_));
 sky130_fd_sc_hd__clkbuf_4 _11905_ (.A(_05754_),
    .X(_05755_));
 sky130_fd_sc_hd__mux2_1 _11906_ (.A0(_05748_),
    .A1(_05753_),
    .S(_05755_),
    .X(_05756_));
 sky130_fd_sc_hd__nand2_1 _11907_ (.A(_05756_),
    .B(_05743_),
    .Y(_05757_));
 sky130_fd_sc_hd__o211a_1 _11908_ (.A1(\result_reg_Lshift[1] ),
    .A2(_05743_),
    .B1(_05672_),
    .C1(_05757_),
    .X(_00309_));
 sky130_fd_sc_hd__a22o_1 _11909_ (.A1(_01158_),
    .A2(_02719_),
    .B1(_02730_),
    .B2(_05749_),
    .X(_05758_));
 sky130_fd_sc_hd__a21o_2 _11910_ (.A1(_05744_),
    .A2(_02711_),
    .B1(_05758_),
    .X(_05759_));
 sky130_fd_sc_hd__nand2_1 _11911_ (.A(_02866_),
    .B(_02869_),
    .Y(_05760_));
 sky130_fd_sc_hd__a22o_1 _11912_ (.A1(_01158_),
    .A2(_02881_),
    .B1(_02891_),
    .B2(_05749_),
    .X(_05761_));
 sky130_fd_sc_hd__a21o_2 _11913_ (.A1(_05744_),
    .A2(_05760_),
    .B1(_05761_),
    .X(_05762_));
 sky130_fd_sc_hd__mux2_1 _11914_ (.A0(_05759_),
    .A1(_05762_),
    .S(_05755_),
    .X(_05763_));
 sky130_fd_sc_hd__nand2_1 _11915_ (.A(_05763_),
    .B(_05743_),
    .Y(_05764_));
 sky130_fd_sc_hd__o211a_1 _11916_ (.A1(\result_reg_Lshift[2] ),
    .A2(_05743_),
    .B1(_05672_),
    .C1(_05764_),
    .X(_00310_));
 sky130_fd_sc_hd__nand2_1 _11917_ (.A(_00591_),
    .B(_05754_),
    .Y(_05765_));
 sky130_fd_sc_hd__buf_4 _11918_ (.A(_05749_),
    .X(_05766_));
 sky130_fd_sc_hd__inv_2 _11919_ (.A(_03162_),
    .Y(_05767_));
 sky130_fd_sc_hd__nor2_1 _11920_ (.A(_00591_),
    .B(_05767_),
    .Y(_05768_));
 sky130_fd_sc_hd__a221o_2 _11921_ (.A1(_05745_),
    .A2(_03169_),
    .B1(_03155_),
    .B2(_05766_),
    .C1(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__o22a_1 _11922_ (.A1(_05755_),
    .A2(_05753_),
    .B1(_05765_),
    .B2(_05769_),
    .X(_05770_));
 sky130_fd_sc_hd__clkbuf_4 _11923_ (.A(_05741_),
    .X(_05771_));
 sky130_fd_sc_hd__nor2_1 _11924_ (.A(\result_reg_Lshift[3] ),
    .B(_05771_),
    .Y(_05772_));
 sky130_fd_sc_hd__a211o_1 _11925_ (.A1(_05770_),
    .A2(_05771_),
    .B1(_05710_),
    .C1(_05772_),
    .X(_05773_));
 sky130_fd_sc_hd__inv_2 _11926_ (.A(_05773_),
    .Y(_00311_));
 sky130_fd_sc_hd__inv_2 _11927_ (.A(_05741_),
    .Y(_05774_));
 sky130_fd_sc_hd__buf_4 _11928_ (.A(_00635_),
    .X(_05775_));
 sky130_fd_sc_hd__nand2_1 _11929_ (.A(_00591_),
    .B(_02118_),
    .Y(_05776_));
 sky130_fd_sc_hd__inv_2 _11930_ (.A(_03128_),
    .Y(_05777_));
 sky130_fd_sc_hd__nor2_1 _11931_ (.A(_00591_),
    .B(_05777_),
    .Y(_05778_));
 sky130_fd_sc_hd__a221o_2 _11932_ (.A1(_03122_),
    .A2(_05745_),
    .B1(_03141_),
    .B2(_05749_),
    .C1(_05778_),
    .X(_05779_));
 sky130_fd_sc_hd__o22ai_2 _11933_ (.A1(_05762_),
    .A2(_05776_),
    .B1(_02118_),
    .B2(_05779_),
    .Y(_05780_));
 sky130_fd_sc_hd__nor2_1 _11934_ (.A(_05774_),
    .B(_05780_),
    .Y(_05781_));
 sky130_fd_sc_hd__a211o_1 _11935_ (.A1(_00806_),
    .A2(_05774_),
    .B1(_05775_),
    .C1(_05781_),
    .X(_05782_));
 sky130_fd_sc_hd__inv_2 _11936_ (.A(_05782_),
    .Y(_00312_));
 sky130_fd_sc_hd__nand2_1 _11937_ (.A(_03082_),
    .B(_03084_),
    .Y(_05783_));
 sky130_fd_sc_hd__a22o_1 _11938_ (.A1(_01158_),
    .A2(_03091_),
    .B1(_03102_),
    .B2(_05749_),
    .X(_05784_));
 sky130_fd_sc_hd__a21o_2 _11939_ (.A1(_05744_),
    .A2(_05783_),
    .B1(_05784_),
    .X(_05785_));
 sky130_fd_sc_hd__mux2_1 _11940_ (.A0(_05769_),
    .A1(_05785_),
    .S(_05755_),
    .X(_05786_));
 sky130_fd_sc_hd__nand2_1 _11941_ (.A(_05786_),
    .B(_05771_),
    .Y(_05787_));
 sky130_fd_sc_hd__o211a_1 _11942_ (.A1(\result_reg_Lshift[5] ),
    .A2(_05743_),
    .B1(_05672_),
    .C1(_05787_),
    .X(_00313_));
 sky130_fd_sc_hd__nand2_1 _11943_ (.A(_03072_),
    .B(_05749_),
    .Y(_05788_));
 sky130_fd_sc_hd__nand2_1 _11944_ (.A(_03054_),
    .B(_03056_),
    .Y(_05789_));
 sky130_fd_sc_hd__nand2_1 _11945_ (.A(_05789_),
    .B(_00590_),
    .Y(_05790_));
 sky130_fd_sc_hd__nand2_1 _11946_ (.A(_03063_),
    .B(_01158_),
    .Y(_05791_));
 sky130_fd_sc_hd__and3_2 _11947_ (.A(_05788_),
    .B(_05790_),
    .C(_05791_),
    .X(_05792_));
 sky130_fd_sc_hd__inv_2 _11948_ (.A(_05792_),
    .Y(_05793_));
 sky130_fd_sc_hd__mux2_1 _11949_ (.A0(_05779_),
    .A1(_05793_),
    .S(_05755_),
    .X(_05794_));
 sky130_fd_sc_hd__nand2_1 _11950_ (.A(_05794_),
    .B(_05771_),
    .Y(_05795_));
 sky130_fd_sc_hd__o211a_1 _11951_ (.A1(\result_reg_Lshift[6] ),
    .A2(_05743_),
    .B1(_05672_),
    .C1(_05795_),
    .X(_00314_));
 sky130_fd_sc_hd__nand2_1 _11952_ (.A(_03824_),
    .B(_01158_),
    .Y(_05796_));
 sky130_fd_sc_hd__nand2_1 _11953_ (.A(_03819_),
    .B(_00590_),
    .Y(_05797_));
 sky130_fd_sc_hd__nand2_1 _11954_ (.A(_03831_),
    .B(_00589_),
    .Y(_05798_));
 sky130_fd_sc_hd__and3_1 _11955_ (.A(_05796_),
    .B(_05797_),
    .C(_05798_),
    .X(_05799_));
 sky130_fd_sc_hd__nor2_1 _11956_ (.A(_05755_),
    .B(_05785_),
    .Y(_05800_));
 sky130_fd_sc_hd__a31o_1 _11957_ (.A1(_05799_),
    .A2(_05766_),
    .A3(_05755_),
    .B1(_05800_),
    .X(_05801_));
 sky130_fd_sc_hd__nand2_1 _11958_ (.A(_05774_),
    .B(_00901_),
    .Y(_05802_));
 sky130_fd_sc_hd__o211a_1 _11959_ (.A1(_05774_),
    .A2(_05801_),
    .B1(_05672_),
    .C1(_05802_),
    .X(_00315_));
 sky130_fd_sc_hd__inv_2 _11960_ (.A(_03854_),
    .Y(_05803_));
 sky130_fd_sc_hd__nor2_1 _11961_ (.A(_01554_),
    .B(_05803_),
    .Y(_05804_));
 sky130_fd_sc_hd__a221o_2 _11962_ (.A1(_03840_),
    .A2(_05744_),
    .B1(_03846_),
    .B2(_05745_),
    .C1(_05804_),
    .X(_05805_));
 sky130_fd_sc_hd__nor2_1 _11963_ (.A(_02118_),
    .B(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__a31o_1 _11964_ (.A1(_05766_),
    .A2(_02118_),
    .A3(_05792_),
    .B1(_05806_),
    .X(_05807_));
 sky130_fd_sc_hd__clkbuf_4 _11965_ (.A(_01148_),
    .X(_05808_));
 sky130_fd_sc_hd__nand2_1 _11966_ (.A(_05774_),
    .B(_00923_),
    .Y(_05809_));
 sky130_fd_sc_hd__o211a_1 _11967_ (.A1(_05774_),
    .A2(_05807_),
    .B1(_05808_),
    .C1(_05809_),
    .X(_00316_));
 sky130_fd_sc_hd__nor2_1 _11968_ (.A(_01554_),
    .B(_03874_),
    .Y(_05810_));
 sky130_fd_sc_hd__a221oi_4 _11969_ (.A1(_00590_),
    .A2(_04552_),
    .B1(_04546_),
    .B2(_01158_),
    .C1(_05810_),
    .Y(_05811_));
 sky130_fd_sc_hd__inv_2 _11970_ (.A(_05811_),
    .Y(_05812_));
 sky130_fd_sc_hd__inv_2 _11971_ (.A(_05799_),
    .Y(_05813_));
 sky130_fd_sc_hd__mux2_1 _11972_ (.A0(_05812_),
    .A1(_05813_),
    .S(_02118_),
    .X(_05814_));
 sky130_fd_sc_hd__nand2_1 _11973_ (.A(_05814_),
    .B(_05771_),
    .Y(_05815_));
 sky130_fd_sc_hd__o211a_1 _11974_ (.A1(\result_reg_Lshift[9] ),
    .A2(_05743_),
    .B1(_05808_),
    .C1(_05815_),
    .X(_00317_));
 sky130_fd_sc_hd__nor2_1 _11975_ (.A(_01554_),
    .B(_03866_),
    .Y(_05816_));
 sky130_fd_sc_hd__a221o_2 _11976_ (.A1(_00590_),
    .A2(_04741_),
    .B1(_04735_),
    .B2(_01158_),
    .C1(_05816_),
    .X(_05817_));
 sky130_fd_sc_hd__mux2_1 _11977_ (.A0(_05805_),
    .A1(_05817_),
    .S(_05755_),
    .X(_05818_));
 sky130_fd_sc_hd__nand2_1 _11978_ (.A(_05818_),
    .B(_05771_),
    .Y(_05819_));
 sky130_fd_sc_hd__o211a_1 _11979_ (.A1(\result_reg_Lshift[10] ),
    .A2(_05743_),
    .B1(_05808_),
    .C1(_05819_),
    .X(_00318_));
 sky130_fd_sc_hd__nor2_1 _11980_ (.A(_02139_),
    .B(_04886_),
    .Y(_05820_));
 sky130_fd_sc_hd__a221o_2 _11981_ (.A1(_04891_),
    .A2(_05744_),
    .B1(_04107_),
    .B2(_05766_),
    .C1(_05820_),
    .X(_05821_));
 sky130_fd_sc_hd__o22a_1 _11982_ (.A1(_05755_),
    .A2(_05812_),
    .B1(_05765_),
    .B2(_05821_),
    .X(_05822_));
 sky130_fd_sc_hd__nor2_1 _11983_ (.A(\result_reg_Lshift[11] ),
    .B(_05741_),
    .Y(_05823_));
 sky130_fd_sc_hd__a211o_1 _11984_ (.A1(_05822_),
    .A2(_05771_),
    .B1(_05775_),
    .C1(_05823_),
    .X(_05824_));
 sky130_fd_sc_hd__inv_2 _11985_ (.A(_05824_),
    .Y(_00319_));
 sky130_fd_sc_hd__inv_2 _11986_ (.A(_04969_),
    .Y(_05825_));
 sky130_fd_sc_hd__nor2_1 _11987_ (.A(_01162_),
    .B(_05825_),
    .Y(_05826_));
 sky130_fd_sc_hd__a221oi_2 _11988_ (.A1(_04963_),
    .A2(_00590_),
    .B1(_04047_),
    .B2(_05749_),
    .C1(_05826_),
    .Y(_05827_));
 sky130_fd_sc_hd__inv_2 _11989_ (.A(_05827_),
    .Y(_05828_));
 sky130_fd_sc_hd__o22a_1 _11990_ (.A1(_05776_),
    .A2(_05817_),
    .B1(_02118_),
    .B2(_05828_),
    .X(_05829_));
 sky130_fd_sc_hd__nor2_1 _11991_ (.A(\result_reg_Lshift[12] ),
    .B(_05741_),
    .Y(_05830_));
 sky130_fd_sc_hd__a211o_1 _11992_ (.A1(_05829_),
    .A2(_05771_),
    .B1(_05775_),
    .C1(_05830_),
    .X(_05831_));
 sky130_fd_sc_hd__inv_2 _11993_ (.A(_05831_),
    .Y(_00320_));
 sky130_fd_sc_hd__and2_1 _11994_ (.A(_04058_),
    .B(_00590_),
    .X(_05832_));
 sky130_fd_sc_hd__a221o_2 _11995_ (.A1(_04071_),
    .A2(_05749_),
    .B1(_04064_),
    .B2(_05745_),
    .C1(_05832_),
    .X(_05833_));
 sky130_fd_sc_hd__mux2_1 _11996_ (.A0(_05821_),
    .A1(_05833_),
    .S(_05754_),
    .X(_05834_));
 sky130_fd_sc_hd__nand2_1 _11997_ (.A(_05834_),
    .B(_05771_),
    .Y(_05835_));
 sky130_fd_sc_hd__o211a_1 _11998_ (.A1(\result_reg_Lshift[13] ),
    .A2(_05743_),
    .B1(_05808_),
    .C1(_05835_),
    .X(_00321_));
 sky130_fd_sc_hd__and2_1 _11999_ (.A(_04078_),
    .B(_04080_),
    .X(_05836_));
 sky130_fd_sc_hd__nor2_1 _12000_ (.A(_00591_),
    .B(_05836_),
    .Y(_05837_));
 sky130_fd_sc_hd__a221o_1 _12001_ (.A1(_04093_),
    .A2(_05749_),
    .B1(_04086_),
    .B2(_05745_),
    .C1(_05837_),
    .X(_05838_));
 sky130_fd_sc_hd__mux2_1 _12002_ (.A0(_05828_),
    .A1(_05838_),
    .S(_05754_),
    .X(_05839_));
 sky130_fd_sc_hd__nand2_1 _12003_ (.A(_05839_),
    .B(_05771_),
    .Y(_05840_));
 sky130_fd_sc_hd__o211a_1 _12004_ (.A1(\result_reg_Lshift[14] ),
    .A2(_05743_),
    .B1(_05808_),
    .C1(_05840_),
    .X(_00322_));
 sky130_fd_sc_hd__nor2_1 _12005_ (.A(_05755_),
    .B(_05833_),
    .Y(_05841_));
 sky130_fd_sc_hd__nand2_1 _12006_ (.A(_05774_),
    .B(_01103_),
    .Y(_05842_));
 sky130_fd_sc_hd__o211a_1 _12007_ (.A1(_05774_),
    .A2(_05841_),
    .B1(_05808_),
    .C1(_05842_),
    .X(_00323_));
 sky130_fd_sc_hd__nand2_2 _12008_ (.A(_00640_),
    .B(_05667_),
    .Y(_05843_));
 sky130_fd_sc_hd__clkbuf_4 _12009_ (.A(_05843_),
    .X(_05844_));
 sky130_fd_sc_hd__nor2_1 _12010_ (.A(_02118_),
    .B(_05759_),
    .Y(_05845_));
 sky130_fd_sc_hd__nand2_1 _12011_ (.A(_05844_),
    .B(_00658_),
    .Y(_05846_));
 sky130_fd_sc_hd__o211a_1 _12012_ (.A1(_05844_),
    .A2(_05845_),
    .B1(_05808_),
    .C1(_05846_),
    .X(_00324_));
 sky130_fd_sc_hd__inv_2 _12013_ (.A(_05843_),
    .Y(_05847_));
 sky130_fd_sc_hd__buf_2 _12014_ (.A(_05847_),
    .X(_05848_));
 sky130_fd_sc_hd__nand2_1 _12015_ (.A(_05756_),
    .B(_05848_),
    .Y(_05849_));
 sky130_fd_sc_hd__o211a_1 _12016_ (.A1(\result_reg_Rshift[1] ),
    .A2(_05848_),
    .B1(_05808_),
    .C1(_05849_),
    .X(_00325_));
 sky130_fd_sc_hd__nand2_1 _12017_ (.A(_05763_),
    .B(_05848_),
    .Y(_05850_));
 sky130_fd_sc_hd__o211a_1 _12018_ (.A1(\result_reg_Rshift[2] ),
    .A2(_05848_),
    .B1(_05808_),
    .C1(_05850_),
    .X(_00326_));
 sky130_fd_sc_hd__clkbuf_4 _12019_ (.A(_05847_),
    .X(_05851_));
 sky130_fd_sc_hd__nor2_1 _12020_ (.A(\result_reg_Rshift[3] ),
    .B(_05851_),
    .Y(_05852_));
 sky130_fd_sc_hd__a211o_1 _12021_ (.A1(_05770_),
    .A2(_05851_),
    .B1(_05775_),
    .C1(_05852_),
    .X(_05853_));
 sky130_fd_sc_hd__inv_2 _12022_ (.A(_05853_),
    .Y(_00327_));
 sky130_fd_sc_hd__nor2_1 _12023_ (.A(_05844_),
    .B(_05780_),
    .Y(_05854_));
 sky130_fd_sc_hd__a211o_1 _12024_ (.A1(_00805_),
    .A2(_05844_),
    .B1(_05775_),
    .C1(_05854_),
    .X(_05855_));
 sky130_fd_sc_hd__inv_2 _12025_ (.A(_05855_),
    .Y(_00328_));
 sky130_fd_sc_hd__nand2_1 _12026_ (.A(_05786_),
    .B(_05851_),
    .Y(_05856_));
 sky130_fd_sc_hd__o211a_1 _12027_ (.A1(\result_reg_Rshift[5] ),
    .A2(_05848_),
    .B1(_05808_),
    .C1(_05856_),
    .X(_00329_));
 sky130_fd_sc_hd__clkbuf_4 _12028_ (.A(_01148_),
    .X(_05857_));
 sky130_fd_sc_hd__nand2_1 _12029_ (.A(_05794_),
    .B(_05851_),
    .Y(_05858_));
 sky130_fd_sc_hd__o211a_1 _12030_ (.A1(\result_reg_Rshift[6] ),
    .A2(_05848_),
    .B1(_05857_),
    .C1(_05858_),
    .X(_00330_));
 sky130_fd_sc_hd__nand2_1 _12031_ (.A(_05844_),
    .B(_00900_),
    .Y(_05859_));
 sky130_fd_sc_hd__o211a_1 _12032_ (.A1(_05844_),
    .A2(_05801_),
    .B1(_05857_),
    .C1(_05859_),
    .X(_00331_));
 sky130_fd_sc_hd__nand2_1 _12033_ (.A(_05844_),
    .B(_00922_),
    .Y(_05860_));
 sky130_fd_sc_hd__o211a_1 _12034_ (.A1(_05844_),
    .A2(_05807_),
    .B1(_05857_),
    .C1(_05860_),
    .X(_00332_));
 sky130_fd_sc_hd__nand2_1 _12035_ (.A(_05814_),
    .B(_05851_),
    .Y(_05861_));
 sky130_fd_sc_hd__o211a_1 _12036_ (.A1(\result_reg_Rshift[9] ),
    .A2(_05848_),
    .B1(_05857_),
    .C1(_05861_),
    .X(_00333_));
 sky130_fd_sc_hd__nand2_1 _12037_ (.A(_05818_),
    .B(_05851_),
    .Y(_05862_));
 sky130_fd_sc_hd__o211a_1 _12038_ (.A1(\result_reg_Rshift[10] ),
    .A2(_05848_),
    .B1(_05857_),
    .C1(_05862_),
    .X(_00334_));
 sky130_fd_sc_hd__nor2_1 _12039_ (.A(\result_reg_Rshift[11] ),
    .B(_05847_),
    .Y(_05863_));
 sky130_fd_sc_hd__a211o_1 _12040_ (.A1(_05822_),
    .A2(_05851_),
    .B1(_05775_),
    .C1(_05863_),
    .X(_05864_));
 sky130_fd_sc_hd__inv_2 _12041_ (.A(_05864_),
    .Y(_00335_));
 sky130_fd_sc_hd__nor2_1 _12042_ (.A(\result_reg_Rshift[12] ),
    .B(_05847_),
    .Y(_05865_));
 sky130_fd_sc_hd__a211o_1 _12043_ (.A1(_05829_),
    .A2(_05851_),
    .B1(_05775_),
    .C1(_05865_),
    .X(_05866_));
 sky130_fd_sc_hd__inv_2 _12044_ (.A(_05866_),
    .Y(_00336_));
 sky130_fd_sc_hd__nand2_1 _12045_ (.A(_05834_),
    .B(_05851_),
    .Y(_05867_));
 sky130_fd_sc_hd__o211a_1 _12046_ (.A1(\result_reg_Rshift[13] ),
    .A2(_05848_),
    .B1(_05857_),
    .C1(_05867_),
    .X(_00337_));
 sky130_fd_sc_hd__nand2_1 _12047_ (.A(_05839_),
    .B(_05851_),
    .Y(_05868_));
 sky130_fd_sc_hd__o211a_1 _12048_ (.A1(\result_reg_Rshift[14] ),
    .A2(_05848_),
    .B1(_05857_),
    .C1(_05868_),
    .X(_00338_));
 sky130_fd_sc_hd__nand2_1 _12049_ (.A(_05844_),
    .B(_01102_),
    .Y(_05869_));
 sky130_fd_sc_hd__o211a_1 _12050_ (.A1(_05844_),
    .A2(_05841_),
    .B1(_05857_),
    .C1(_05869_),
    .X(_00339_));
 sky130_fd_sc_hd__nor2_1 _12051_ (.A(_00639_),
    .B(_00572_),
    .Y(_05870_));
 sky130_fd_sc_hd__and3_2 _12052_ (.A(_05870_),
    .B(_00555_),
    .C(_05667_),
    .X(_05871_));
 sky130_fd_sc_hd__inv_2 _12053_ (.A(_05871_),
    .Y(_05872_));
 sky130_fd_sc_hd__clkbuf_4 _12054_ (.A(_05872_),
    .X(_05873_));
 sky130_fd_sc_hd__and3_1 _12055_ (.A(_02613_),
    .B(_02615_),
    .C(_01666_),
    .X(_05874_));
 sky130_fd_sc_hd__nand2_1 _12056_ (.A(_05874_),
    .B(_05746_),
    .Y(_05875_));
 sky130_fd_sc_hd__nand2_1 _12057_ (.A(_02601_),
    .B(_02604_),
    .Y(_05876_));
 sky130_fd_sc_hd__or3_1 _12058_ (.A(_01200_),
    .B(_05876_),
    .C(_02550_),
    .X(_05877_));
 sky130_fd_sc_hd__clkbuf_4 _12059_ (.A(_05871_),
    .X(_05878_));
 sky130_fd_sc_hd__or3_1 _12060_ (.A(_00525_),
    .B(_02538_),
    .C(_02595_),
    .X(_05879_));
 sky130_fd_sc_hd__and4_1 _12061_ (.A(_05875_),
    .B(_05877_),
    .C(_05878_),
    .D(_05879_),
    .X(_05880_));
 sky130_fd_sc_hd__a211oi_1 _12062_ (.A1(_01209_),
    .A2(_05873_),
    .B1(_05775_),
    .C1(_05880_),
    .Y(_00340_));
 sky130_fd_sc_hd__clkbuf_4 _12063_ (.A(_01200_),
    .X(_05881_));
 sky130_fd_sc_hd__nand2_1 _12064_ (.A(_02667_),
    .B(_02670_),
    .Y(_05882_));
 sky130_fd_sc_hd__or3_1 _12065_ (.A(_05881_),
    .B(_05882_),
    .C(_02719_),
    .X(_05883_));
 sky130_fd_sc_hd__nor2_1 _12066_ (.A(_01578_),
    .B(_02730_),
    .Y(_05884_));
 sky130_fd_sc_hd__nand2_1 _12067_ (.A(_05884_),
    .B(_02682_),
    .Y(_05885_));
 sky130_fd_sc_hd__or3_1 _12068_ (.A(_00525_),
    .B(_02711_),
    .C(_02661_),
    .X(_05886_));
 sky130_fd_sc_hd__and4_1 _12069_ (.A(_05883_),
    .B(_05885_),
    .C(_05886_),
    .D(_05878_),
    .X(_05887_));
 sky130_fd_sc_hd__a211oi_1 _12070_ (.A1(_00715_),
    .A2(_05873_),
    .B1(_05775_),
    .C1(_05887_),
    .Y(_00341_));
 sky130_fd_sc_hd__clkbuf_4 _12071_ (.A(_01578_),
    .X(_05888_));
 sky130_fd_sc_hd__nand2_1 _12072_ (.A(_02766_),
    .B(_02769_),
    .Y(_05889_));
 sky130_fd_sc_hd__or3_1 _12073_ (.A(_01200_),
    .B(_05889_),
    .C(_02807_),
    .X(_05890_));
 sky130_fd_sc_hd__o31a_1 _12074_ (.A1(_05888_),
    .A2(_02817_),
    .A3(_02781_),
    .B1(_05890_),
    .X(_05891_));
 sky130_fd_sc_hd__clkbuf_4 _12075_ (.A(_00525_),
    .X(_05892_));
 sky130_fd_sc_hd__o31a_1 _12076_ (.A1(_05892_),
    .A2(_05750_),
    .A3(_02760_),
    .B1(_05878_),
    .X(_05893_));
 sky130_fd_sc_hd__a221oi_1 _12077_ (.A1(_01282_),
    .A2(_05873_),
    .B1(_05891_),
    .B2(_05893_),
    .C1(_02650_),
    .Y(_00342_));
 sky130_fd_sc_hd__clkbuf_4 _12078_ (.A(_05878_),
    .X(_05894_));
 sky130_fd_sc_hd__or3_1 _12079_ (.A(_05881_),
    .B(_02923_),
    .C(_02881_),
    .X(_05895_));
 sky130_fd_sc_hd__nand2_1 _12080_ (.A(_05895_),
    .B(_05894_),
    .Y(_05896_));
 sky130_fd_sc_hd__or3_1 _12081_ (.A(_05892_),
    .B(_02933_),
    .C(_05760_),
    .X(_05897_));
 sky130_fd_sc_hd__nor2_1 _12082_ (.A(_05888_),
    .B(_02891_),
    .Y(_05898_));
 sky130_fd_sc_hd__nand2_1 _12083_ (.A(_02944_),
    .B(_05898_),
    .Y(_05899_));
 sky130_fd_sc_hd__nand2_1 _12084_ (.A(_05897_),
    .B(_05899_),
    .Y(_05900_));
 sky130_fd_sc_hd__o221a_1 _12085_ (.A1(\result_reg_and[3] ),
    .A2(_05894_),
    .B1(_05896_),
    .B2(_05900_),
    .C1(_02125_),
    .X(_00343_));
 sky130_fd_sc_hd__a41o_1 _12086_ (.A1(_05767_),
    .A2(_00524_),
    .A3(_02994_),
    .A4(_02997_),
    .B1(_05872_),
    .X(_05901_));
 sky130_fd_sc_hd__inv_2 _12087_ (.A(_03169_),
    .Y(_05902_));
 sky130_fd_sc_hd__and2_1 _12088_ (.A(_03003_),
    .B(_03006_),
    .X(_05903_));
 sky130_fd_sc_hd__buf_4 _12089_ (.A(_01666_),
    .X(_05904_));
 sky130_fd_sc_hd__nor2_1 _12090_ (.A(_03015_),
    .B(_03155_),
    .Y(_05905_));
 sky130_fd_sc_hd__a32o_1 _12091_ (.A1(_05902_),
    .A2(_01243_),
    .A3(_05903_),
    .B1(_05904_),
    .B2(_05905_),
    .X(_05906_));
 sky130_fd_sc_hd__o221a_1 _12092_ (.A1(\result_reg_and[4] ),
    .A2(_05894_),
    .B1(_05901_),
    .B2(_05906_),
    .C1(_02125_),
    .X(_00344_));
 sky130_fd_sc_hd__clkbuf_4 _12093_ (.A(_05892_),
    .X(_05907_));
 sky130_fd_sc_hd__o31ai_1 _12094_ (.A1(_05907_),
    .A2(_03328_),
    .A3(_03128_),
    .B1(_05894_),
    .Y(_05908_));
 sky130_fd_sc_hd__and2_1 _12095_ (.A(_03333_),
    .B(_03335_),
    .X(_05909_));
 sky130_fd_sc_hd__or3b_1 _12096_ (.A(_05881_),
    .B(_03122_),
    .C_N(_05909_),
    .X(_05910_));
 sky130_fd_sc_hd__o31ai_1 _12097_ (.A1(_05888_),
    .A2(_03141_),
    .A3(_03346_),
    .B1(_05910_),
    .Y(_05911_));
 sky130_fd_sc_hd__o221a_1 _12098_ (.A1(\result_reg_and[5] ),
    .A2(_05894_),
    .B1(_05908_),
    .B2(_05911_),
    .C1(_02125_),
    .X(_00345_));
 sky130_fd_sc_hd__or3_1 _12099_ (.A(_01200_),
    .B(_03482_),
    .C(_03091_),
    .X(_05912_));
 sky130_fd_sc_hd__o31a_1 _12100_ (.A1(_01578_),
    .A2(_03102_),
    .A3(_03502_),
    .B1(_05912_),
    .X(_05913_));
 sky130_fd_sc_hd__o31a_1 _12101_ (.A1(_05892_),
    .A2(_03489_),
    .A3(_05783_),
    .B1(_05878_),
    .X(_05914_));
 sky130_fd_sc_hd__a221oi_1 _12102_ (.A1(_01359_),
    .A2(_05873_),
    .B1(_05913_),
    .B2(_05914_),
    .C1(_02650_),
    .Y(_00346_));
 sky130_fd_sc_hd__or3_1 _12103_ (.A(_01578_),
    .B(_03072_),
    .C(_03647_),
    .X(_05915_));
 sky130_fd_sc_hd__or3_1 _12104_ (.A(_01200_),
    .B(_03063_),
    .C(_03632_),
    .X(_05916_));
 sky130_fd_sc_hd__or3_1 _12105_ (.A(_00525_),
    .B(_03639_),
    .C(_05789_),
    .X(_05917_));
 sky130_fd_sc_hd__and4_1 _12106_ (.A(_05915_),
    .B(_05878_),
    .C(_05916_),
    .D(_05917_),
    .X(_05918_));
 sky130_fd_sc_hd__a211oi_1 _12107_ (.A1(_01776_),
    .A2(_05873_),
    .B1(_02115_),
    .C1(_05918_),
    .Y(_00347_));
 sky130_fd_sc_hd__or3_1 _12108_ (.A(_05892_),
    .B(_03780_),
    .C(_03819_),
    .X(_05919_));
 sky130_fd_sc_hd__o31ai_1 _12109_ (.A1(_05888_),
    .A2(_03767_),
    .A3(_03831_),
    .B1(_05919_),
    .Y(_05920_));
 sky130_fd_sc_hd__o31ai_1 _12110_ (.A1(_05881_),
    .A2(_03824_),
    .A3(_03775_),
    .B1(_05894_),
    .Y(_05921_));
 sky130_fd_sc_hd__o221a_1 _12111_ (.A1(\result_reg_and[8] ),
    .A2(_05894_),
    .B1(_05920_),
    .B2(_05921_),
    .C1(_02125_),
    .X(_00348_));
 sky130_fd_sc_hd__nor2_1 _12112_ (.A(_01578_),
    .B(_04305_),
    .Y(_05922_));
 sky130_fd_sc_hd__nand2_1 _12113_ (.A(_05922_),
    .B(_05803_),
    .Y(_05923_));
 sky130_fd_sc_hd__or3_1 _12114_ (.A(_01200_),
    .B(_04288_),
    .C(_03846_),
    .X(_05924_));
 sky130_fd_sc_hd__or3_1 _12115_ (.A(_00525_),
    .B(_03840_),
    .C(_04294_),
    .X(_05925_));
 sky130_fd_sc_hd__and4_1 _12116_ (.A(_05923_),
    .B(_05924_),
    .C(_05925_),
    .D(_05871_),
    .X(_05926_));
 sky130_fd_sc_hd__a211oi_1 _12117_ (.A1(_01407_),
    .A2(_05873_),
    .B1(_02115_),
    .C1(_05926_),
    .Y(_00349_));
 sky130_fd_sc_hd__or3_1 _12118_ (.A(_01200_),
    .B(_04483_),
    .C(_04546_),
    .X(_05927_));
 sky130_fd_sc_hd__nor2_1 _12119_ (.A(_01578_),
    .B(_04490_),
    .Y(_05928_));
 sky130_fd_sc_hd__nand2_1 _12120_ (.A(_05928_),
    .B(_03874_),
    .Y(_05929_));
 sky130_fd_sc_hd__or3_1 _12121_ (.A(_00525_),
    .B(_04552_),
    .C(_04477_),
    .X(_05930_));
 sky130_fd_sc_hd__and4_1 _12122_ (.A(_05927_),
    .B(_05929_),
    .C(_05930_),
    .D(_05871_),
    .X(_05931_));
 sky130_fd_sc_hd__a211oi_1 _12123_ (.A1(_01831_),
    .A2(_05873_),
    .B1(_02115_),
    .C1(_05931_),
    .Y(_00350_));
 sky130_fd_sc_hd__nand2_1 _12124_ (.A(_04671_),
    .B(_03866_),
    .Y(_05932_));
 sky130_fd_sc_hd__or3_1 _12125_ (.A(_00525_),
    .B(_04741_),
    .C(_04677_),
    .X(_05933_));
 sky130_fd_sc_hd__or3_1 _12126_ (.A(_05881_),
    .B(_04683_),
    .C(_04735_),
    .X(_05934_));
 sky130_fd_sc_hd__o2111a_1 _12127_ (.A1(_05888_),
    .A2(_05932_),
    .B1(_05878_),
    .C1(_05933_),
    .D1(_05934_),
    .X(_05935_));
 sky130_fd_sc_hd__a211oi_1 _12128_ (.A1(_01851_),
    .A2(_05873_),
    .B1(_02115_),
    .C1(_05935_),
    .Y(_00351_));
 sky130_fd_sc_hd__o31ai_1 _12129_ (.A1(_05907_),
    .A2(_04847_),
    .A3(_04891_),
    .B1(_05878_),
    .Y(_05936_));
 sky130_fd_sc_hd__clkbuf_4 _12130_ (.A(_01243_),
    .X(_05937_));
 sky130_fd_sc_hd__nor2_1 _12131_ (.A(_01578_),
    .B(_04107_),
    .Y(_05938_));
 sky130_fd_sc_hd__a32o_1 _12132_ (.A1(_05937_),
    .A2(_04886_),
    .A3(_04842_),
    .B1(_05938_),
    .B2(_04836_),
    .X(_05939_));
 sky130_fd_sc_hd__clkbuf_4 _12133_ (.A(_05682_),
    .X(_05940_));
 sky130_fd_sc_hd__o221a_1 _12134_ (.A1(\result_reg_and[12] ),
    .A2(_05894_),
    .B1(_05936_),
    .B2(_05939_),
    .C1(_05940_),
    .X(_00352_));
 sky130_fd_sc_hd__o31ai_1 _12135_ (.A1(_05907_),
    .A2(_04963_),
    .A3(_05147_),
    .B1(_05878_),
    .Y(_05941_));
 sky130_fd_sc_hd__nor2_1 _12136_ (.A(_05881_),
    .B(_05141_),
    .Y(_05942_));
 sky130_fd_sc_hd__nor2_1 _12137_ (.A(_05888_),
    .B(_04047_),
    .Y(_05943_));
 sky130_fd_sc_hd__a22o_1 _12138_ (.A1(_05825_),
    .A2(_05942_),
    .B1(_05943_),
    .B2(_05154_),
    .X(_05944_));
 sky130_fd_sc_hd__o221a_1 _12139_ (.A1(\result_reg_and[13] ),
    .A2(_05894_),
    .B1(_05941_),
    .B2(_05944_),
    .C1(_05940_),
    .X(_00353_));
 sky130_fd_sc_hd__or3_1 _12140_ (.A(_01200_),
    .B(_04064_),
    .C(_05324_),
    .X(_05945_));
 sky130_fd_sc_hd__or3_1 _12141_ (.A(_00525_),
    .B(_04058_),
    .C(_05329_),
    .X(_05946_));
 sky130_fd_sc_hd__nor2_1 _12142_ (.A(_01578_),
    .B(_04071_),
    .Y(_05947_));
 sky130_fd_sc_hd__nand2_1 _12143_ (.A(_05947_),
    .B(_05338_),
    .Y(_05948_));
 sky130_fd_sc_hd__and4_1 _12144_ (.A(_05945_),
    .B(_05946_),
    .C(_05878_),
    .D(_05948_),
    .X(_05949_));
 sky130_fd_sc_hd__a211oi_1 _12145_ (.A1(_01499_),
    .A2(_05873_),
    .B1(_02115_),
    .C1(_05949_),
    .Y(_00354_));
 sky130_fd_sc_hd__a31o_1 _12146_ (.A1(_05506_),
    .A2(_00524_),
    .A3(_05836_),
    .B1(_05873_),
    .X(_05950_));
 sky130_fd_sc_hd__nor2_1 _12147_ (.A(_05888_),
    .B(_04093_),
    .Y(_05951_));
 sky130_fd_sc_hd__nor2_1 _12148_ (.A(_05881_),
    .B(_04086_),
    .Y(_05952_));
 sky130_fd_sc_hd__a22o_1 _12149_ (.A1(_05515_),
    .A2(_05951_),
    .B1(_05499_),
    .B2(_05952_),
    .X(_05953_));
 sky130_fd_sc_hd__o221a_1 _12150_ (.A1(\result_reg_and[15] ),
    .A2(_05894_),
    .B1(_05950_),
    .B2(_05953_),
    .C1(_05940_),
    .X(_00355_));
 sky130_fd_sc_hd__nor2_1 _12151_ (.A(_00554_),
    .B(_05666_),
    .Y(_05954_));
 sky130_fd_sc_hd__inv_2 _12152_ (.A(_05954_),
    .Y(_05955_));
 sky130_fd_sc_hd__or4_1 _12153_ (.A(_00662_),
    .B(_00572_),
    .C(_05955_),
    .D(_02167_),
    .X(_05956_));
 sky130_fd_sc_hd__clkbuf_4 _12154_ (.A(_05956_),
    .X(_05957_));
 sky130_fd_sc_hd__inv_2 _12155_ (.A(_05957_),
    .Y(_05958_));
 sky130_fd_sc_hd__clkbuf_4 _12156_ (.A(_05958_),
    .X(_05959_));
 sky130_fd_sc_hd__buf_2 _12157_ (.A(_05958_),
    .X(_05960_));
 sky130_fd_sc_hd__a21o_1 _12158_ (.A1(_02538_),
    .A2(_02595_),
    .B1(_05907_),
    .X(_05961_));
 sky130_fd_sc_hd__nand2_1 _12159_ (.A(_05960_),
    .B(_05961_),
    .Y(_05962_));
 sky130_fd_sc_hd__nand2_1 _12160_ (.A(_02550_),
    .B(_05876_),
    .Y(_05963_));
 sky130_fd_sc_hd__a221o_1 _12161_ (.A1(_05904_),
    .A2(_05746_),
    .B1(_01243_),
    .B2(_05963_),
    .C1(_05874_),
    .X(_05964_));
 sky130_fd_sc_hd__o221a_1 _12162_ (.A1(\result_reg_or[0] ),
    .A2(_05959_),
    .B1(_05962_),
    .B2(_05964_),
    .C1(_05940_),
    .X(_00356_));
 sky130_fd_sc_hd__nand2_1 _12163_ (.A(_02711_),
    .B(_02661_),
    .Y(_05965_));
 sky130_fd_sc_hd__nand2_1 _12164_ (.A(_02719_),
    .B(_05882_),
    .Y(_05966_));
 sky130_fd_sc_hd__a22o_1 _12165_ (.A1(_00524_),
    .A2(_05965_),
    .B1(_05966_),
    .B2(_05937_),
    .X(_05967_));
 sky130_fd_sc_hd__a211o_1 _12166_ (.A1(_05904_),
    .A2(_02682_),
    .B1(_05884_),
    .C1(_05957_),
    .X(_05968_));
 sky130_fd_sc_hd__o221a_1 _12167_ (.A1(\result_reg_or[1] ),
    .A2(_05959_),
    .B1(_05967_),
    .B2(_05968_),
    .C1(_05940_),
    .X(_00357_));
 sky130_fd_sc_hd__a21oi_1 _12168_ (.A1(_05750_),
    .A2(_02760_),
    .B1(_05907_),
    .Y(_05969_));
 sky130_fd_sc_hd__nand2_1 _12169_ (.A(_02807_),
    .B(_05889_),
    .Y(_05970_));
 sky130_fd_sc_hd__nand2_1 _12170_ (.A(_02781_),
    .B(_02817_),
    .Y(_05971_));
 sky130_fd_sc_hd__a22o_1 _12171_ (.A1(_01243_),
    .A2(_05970_),
    .B1(_05971_),
    .B2(_01666_),
    .X(_05972_));
 sky130_fd_sc_hd__nand2_1 _12172_ (.A(_05957_),
    .B(_00738_),
    .Y(_05973_));
 sky130_fd_sc_hd__o311a_1 _12173_ (.A1(_05969_),
    .A2(_05972_),
    .A3(_05957_),
    .B1(_04827_),
    .C1(_05973_),
    .X(_00358_));
 sky130_fd_sc_hd__nand2_1 _12174_ (.A(_02933_),
    .B(_05760_),
    .Y(_05974_));
 sky130_fd_sc_hd__nand2_1 _12175_ (.A(_02881_),
    .B(_02923_),
    .Y(_05975_));
 sky130_fd_sc_hd__a22o_1 _12176_ (.A1(_05974_),
    .A2(_00524_),
    .B1(_05937_),
    .B2(_05975_),
    .X(_05976_));
 sky130_fd_sc_hd__a211o_1 _12177_ (.A1(_05904_),
    .A2(_02944_),
    .B1(_05898_),
    .C1(_05957_),
    .X(_05977_));
 sky130_fd_sc_hd__o221a_1 _12178_ (.A1(\result_reg_or[3] ),
    .A2(_05959_),
    .B1(_05976_),
    .B2(_05977_),
    .C1(_05940_),
    .X(_00359_));
 sky130_fd_sc_hd__or2_1 _12179_ (.A(_05903_),
    .B(_05902_),
    .X(_05978_));
 sky130_fd_sc_hd__a21oi_1 _12180_ (.A1(_03162_),
    .A2(_02998_),
    .B1(_05892_),
    .Y(_05979_));
 sky130_fd_sc_hd__a21oi_1 _12181_ (.A1(_03155_),
    .A2(_03015_),
    .B1(_05888_),
    .Y(_05980_));
 sky130_fd_sc_hd__a2111o_1 _12182_ (.A1(_05937_),
    .A2(_05978_),
    .B1(_05979_),
    .C1(_05980_),
    .D1(_05957_),
    .X(_05981_));
 sky130_fd_sc_hd__o211a_1 _12183_ (.A1(\result_reg_or[4] ),
    .A2(_05959_),
    .B1(_05857_),
    .C1(_05981_),
    .X(_00360_));
 sky130_fd_sc_hd__a21o_1 _12184_ (.A1(_03128_),
    .A2(_03328_),
    .B1(_05892_),
    .X(_05982_));
 sky130_fd_sc_hd__o221ai_1 _12185_ (.A1(_05881_),
    .A2(_03122_),
    .B1(_05888_),
    .B2(_03141_),
    .C1(_05982_),
    .Y(_05983_));
 sky130_fd_sc_hd__nor2_1 _12186_ (.A(_05888_),
    .B(_03346_),
    .Y(_05984_));
 sky130_fd_sc_hd__a211o_1 _12187_ (.A1(_05937_),
    .A2(_05909_),
    .B1(_05984_),
    .C1(_05957_),
    .X(_05985_));
 sky130_fd_sc_hd__o221a_1 _12188_ (.A1(\result_reg_or[5] ),
    .A2(_05959_),
    .B1(_05983_),
    .B2(_05985_),
    .C1(_05940_),
    .X(_00361_));
 sky130_fd_sc_hd__nand2_1 _12189_ (.A(_03091_),
    .B(_03482_),
    .Y(_05986_));
 sky130_fd_sc_hd__nand2_1 _12190_ (.A(_03502_),
    .B(_03102_),
    .Y(_05987_));
 sky130_fd_sc_hd__a22o_1 _12191_ (.A1(_05937_),
    .A2(_05986_),
    .B1(_05987_),
    .B2(_05904_),
    .X(_05988_));
 sky130_fd_sc_hd__a21o_1 _12192_ (.A1(_05783_),
    .A2(_03489_),
    .B1(_05907_),
    .X(_05989_));
 sky130_fd_sc_hd__nand2_1 _12193_ (.A(_05960_),
    .B(_05989_),
    .Y(_05990_));
 sky130_fd_sc_hd__o221a_1 _12194_ (.A1(\result_reg_or[6] ),
    .A2(_05959_),
    .B1(_05988_),
    .B2(_05990_),
    .C1(_05940_),
    .X(_00362_));
 sky130_fd_sc_hd__a21o_1 _12195_ (.A1(_05789_),
    .A2(_03639_),
    .B1(_05907_),
    .X(_05991_));
 sky130_fd_sc_hd__nand2_1 _12196_ (.A(_05960_),
    .B(_05991_),
    .Y(_05992_));
 sky130_fd_sc_hd__nand2_1 _12197_ (.A(_03063_),
    .B(_03632_),
    .Y(_05993_));
 sky130_fd_sc_hd__nand2_1 _12198_ (.A(_03647_),
    .B(_03072_),
    .Y(_05994_));
 sky130_fd_sc_hd__a22o_1 _12199_ (.A1(_05937_),
    .A2(_05993_),
    .B1(_05994_),
    .B2(_05904_),
    .X(_05995_));
 sky130_fd_sc_hd__o221a_1 _12200_ (.A1(\result_reg_or[7] ),
    .A2(_05959_),
    .B1(_05992_),
    .B2(_05995_),
    .C1(_05940_),
    .X(_00363_));
 sky130_fd_sc_hd__a21o_1 _12201_ (.A1(_03780_),
    .A2(_03819_),
    .B1(_05907_),
    .X(_05996_));
 sky130_fd_sc_hd__nand2_1 _12202_ (.A(_05960_),
    .B(_05996_),
    .Y(_05997_));
 sky130_fd_sc_hd__nand2_1 _12203_ (.A(_03831_),
    .B(_03767_),
    .Y(_05998_));
 sky130_fd_sc_hd__nand2_1 _12204_ (.A(_03775_),
    .B(_03824_),
    .Y(_05999_));
 sky130_fd_sc_hd__a22o_1 _12205_ (.A1(_05904_),
    .A2(_05998_),
    .B1(_05999_),
    .B2(_05937_),
    .X(_06000_));
 sky130_fd_sc_hd__o221a_1 _12206_ (.A1(\result_reg_or[8] ),
    .A2(_05959_),
    .B1(_05997_),
    .B2(_06000_),
    .C1(_05940_),
    .X(_00364_));
 sky130_fd_sc_hd__a21o_1 _12207_ (.A1(_04294_),
    .A2(_03840_),
    .B1(_05907_),
    .X(_06001_));
 sky130_fd_sc_hd__nand2_1 _12208_ (.A(_05960_),
    .B(_06001_),
    .Y(_06002_));
 sky130_fd_sc_hd__nand2_1 _12209_ (.A(_03846_),
    .B(_04288_),
    .Y(_06003_));
 sky130_fd_sc_hd__a221o_1 _12210_ (.A1(_05904_),
    .A2(_05803_),
    .B1(_01243_),
    .B2(_06003_),
    .C1(_05922_),
    .X(_06004_));
 sky130_fd_sc_hd__o221a_1 _12211_ (.A1(\result_reg_or[9] ),
    .A2(_05960_),
    .B1(_06002_),
    .B2(_06004_),
    .C1(_02101_),
    .X(_00365_));
 sky130_fd_sc_hd__a21o_1 _12212_ (.A1(_04552_),
    .A2(_04477_),
    .B1(_05907_),
    .X(_06005_));
 sky130_fd_sc_hd__nand2_1 _12213_ (.A(_05958_),
    .B(_06005_),
    .Y(_06006_));
 sky130_fd_sc_hd__nand2_1 _12214_ (.A(_04546_),
    .B(_04483_),
    .Y(_06007_));
 sky130_fd_sc_hd__a221o_1 _12215_ (.A1(_03874_),
    .A2(_01666_),
    .B1(_06007_),
    .B2(_01243_),
    .C1(_05928_),
    .X(_06008_));
 sky130_fd_sc_hd__o221a_1 _12216_ (.A1(\result_reg_or[10] ),
    .A2(_05960_),
    .B1(_06006_),
    .B2(_06008_),
    .C1(_02101_),
    .X(_00366_));
 sky130_fd_sc_hd__nand2_1 _12217_ (.A(_04735_),
    .B(_04683_),
    .Y(_06009_));
 sky130_fd_sc_hd__a21oi_1 _12218_ (.A1(_04741_),
    .A2(_04677_),
    .B1(_05892_),
    .Y(_06010_));
 sky130_fd_sc_hd__o21a_1 _12219_ (.A1(_03866_),
    .A2(_04671_),
    .B1(_01666_),
    .X(_06011_));
 sky130_fd_sc_hd__a2111o_1 _12220_ (.A1(_05937_),
    .A2(_06009_),
    .B1(_06010_),
    .C1(_06011_),
    .D1(_05957_),
    .X(_06012_));
 sky130_fd_sc_hd__o211a_1 _12221_ (.A1(\result_reg_or[11] ),
    .A2(_05959_),
    .B1(_05857_),
    .C1(_06012_),
    .X(_00367_));
 sky130_fd_sc_hd__clkbuf_4 _12222_ (.A(_01148_),
    .X(_06013_));
 sky130_fd_sc_hd__or2_1 _12223_ (.A(_04886_),
    .B(_04842_),
    .X(_06014_));
 sky130_fd_sc_hd__a21oi_1 _12224_ (.A1(_04891_),
    .A2(_04847_),
    .B1(_05892_),
    .Y(_06015_));
 sky130_fd_sc_hd__a21o_1 _12225_ (.A1(_04836_),
    .A2(_01666_),
    .B1(_05938_),
    .X(_06016_));
 sky130_fd_sc_hd__a2111o_1 _12226_ (.A1(_05937_),
    .A2(_06014_),
    .B1(_06015_),
    .C1(_05957_),
    .D1(_06016_),
    .X(_06017_));
 sky130_fd_sc_hd__o211a_1 _12227_ (.A1(\result_reg_or[12] ),
    .A2(_05959_),
    .B1(_06013_),
    .C1(_06017_),
    .X(_00368_));
 sky130_fd_sc_hd__a21o_1 _12228_ (.A1(_05141_),
    .A2(_04969_),
    .B1(_05881_),
    .X(_06018_));
 sky130_fd_sc_hd__nand2_1 _12229_ (.A(_05958_),
    .B(_06018_),
    .Y(_06019_));
 sky130_fd_sc_hd__nand2_1 _12230_ (.A(_05147_),
    .B(_04963_),
    .Y(_06020_));
 sky130_fd_sc_hd__a221o_1 _12231_ (.A1(_06020_),
    .A2(_00524_),
    .B1(_05154_),
    .B2(_01666_),
    .C1(_05943_),
    .X(_06021_));
 sky130_fd_sc_hd__o221a_1 _12232_ (.A1(\result_reg_or[13] ),
    .A2(_05960_),
    .B1(_06019_),
    .B2(_06021_),
    .C1(_02101_),
    .X(_00369_));
 sky130_fd_sc_hd__a21o_1 _12233_ (.A1(_05329_),
    .A2(_04058_),
    .B1(_05892_),
    .X(_06022_));
 sky130_fd_sc_hd__nand2_1 _12234_ (.A(_05958_),
    .B(_06022_),
    .Y(_06023_));
 sky130_fd_sc_hd__nand2_1 _12235_ (.A(_05324_),
    .B(_04064_),
    .Y(_06024_));
 sky130_fd_sc_hd__a221o_1 _12236_ (.A1(_06024_),
    .A2(_01243_),
    .B1(_05338_),
    .B2(_01666_),
    .C1(_05947_),
    .X(_06025_));
 sky130_fd_sc_hd__o221a_1 _12237_ (.A1(\result_reg_or[14] ),
    .A2(_05960_),
    .B1(_06023_),
    .B2(_06025_),
    .C1(_02101_),
    .X(_00370_));
 sky130_fd_sc_hd__a21o_1 _12238_ (.A1(_05500_),
    .A2(_04086_),
    .B1(_05881_),
    .X(_06026_));
 sky130_fd_sc_hd__nand2_1 _12239_ (.A(_05958_),
    .B(_06026_),
    .Y(_06027_));
 sky130_fd_sc_hd__or2_1 _12240_ (.A(_05836_),
    .B(_05506_),
    .X(_06028_));
 sky130_fd_sc_hd__a221o_1 _12241_ (.A1(_05904_),
    .A2(_05515_),
    .B1(_06028_),
    .B2(_00524_),
    .C1(_05951_),
    .X(_06029_));
 sky130_fd_sc_hd__o221a_1 _12242_ (.A1(\result_reg_or[15] ),
    .A2(_05960_),
    .B1(_06027_),
    .B2(_06029_),
    .C1(_02101_),
    .X(_00371_));
 sky130_fd_sc_hd__or4_2 _12243_ (.A(_02164_),
    .B(_05955_),
    .C(_02098_),
    .D(_00632_),
    .X(_06030_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12244_ (.A(_06030_),
    .X(_06031_));
 sky130_fd_sc_hd__clkbuf_4 _12245_ (.A(_06031_),
    .X(_06032_));
 sky130_fd_sc_hd__buf_2 _12246_ (.A(_06031_),
    .X(_06033_));
 sky130_fd_sc_hd__nand2_1 _12247_ (.A(_06033_),
    .B(_00652_),
    .Y(_06034_));
 sky130_fd_sc_hd__o211a_1 _12248_ (.A1(_06032_),
    .A2(_05748_),
    .B1(_06013_),
    .C1(_06034_),
    .X(_00372_));
 sky130_fd_sc_hd__nand2_1 _12249_ (.A(_06033_),
    .B(_00689_),
    .Y(_06035_));
 sky130_fd_sc_hd__o211a_1 _12250_ (.A1(_06032_),
    .A2(_05759_),
    .B1(_06013_),
    .C1(_06035_),
    .X(_00373_));
 sky130_fd_sc_hd__nand2_1 _12251_ (.A(_06033_),
    .B(_00752_),
    .Y(_06036_));
 sky130_fd_sc_hd__o211a_1 _12252_ (.A1(_06032_),
    .A2(_05753_),
    .B1(_06013_),
    .C1(_06036_),
    .X(_00374_));
 sky130_fd_sc_hd__nand2_1 _12253_ (.A(_06033_),
    .B(_00778_),
    .Y(_06037_));
 sky130_fd_sc_hd__o211a_1 _12254_ (.A1(_05762_),
    .A2(_06033_),
    .B1(_06013_),
    .C1(_06037_),
    .X(_00375_));
 sky130_fd_sc_hd__nand2_1 _12255_ (.A(_06033_),
    .B(_00804_),
    .Y(_06038_));
 sky130_fd_sc_hd__o211a_1 _12256_ (.A1(_06032_),
    .A2(_05769_),
    .B1(_06013_),
    .C1(_06038_),
    .X(_00376_));
 sky130_fd_sc_hd__buf_2 _12257_ (.A(_06031_),
    .X(_06039_));
 sky130_fd_sc_hd__nand2_1 _12258_ (.A(_06033_),
    .B(_00849_),
    .Y(_06040_));
 sky130_fd_sc_hd__o211a_1 _12259_ (.A1(_06039_),
    .A2(_05779_),
    .B1(_06013_),
    .C1(_06040_),
    .X(_00377_));
 sky130_fd_sc_hd__nand2_1 _12260_ (.A(_06033_),
    .B(_00873_),
    .Y(_06041_));
 sky130_fd_sc_hd__o211a_1 _12261_ (.A1(_06039_),
    .A2(_05785_),
    .B1(_06013_),
    .C1(_06041_),
    .X(_00378_));
 sky130_fd_sc_hd__nand2_1 _12262_ (.A(_06033_),
    .B(_00899_),
    .Y(_06042_));
 sky130_fd_sc_hd__o211a_1 _12263_ (.A1(_06039_),
    .A2(_05793_),
    .B1(_06013_),
    .C1(_06042_),
    .X(_00379_));
 sky130_fd_sc_hd__or2b_1 _12264_ (.A(\result_reg_not[8] ),
    .B_N(_06031_),
    .X(_06043_));
 sky130_fd_sc_hd__o211a_1 _12265_ (.A1(_06039_),
    .A2(_05813_),
    .B1(_06013_),
    .C1(_06043_),
    .X(_00380_));
 sky130_fd_sc_hd__clkbuf_4 _12266_ (.A(_01148_),
    .X(_06044_));
 sky130_fd_sc_hd__nand2_1 _12267_ (.A(_06033_),
    .B(_00948_),
    .Y(_06045_));
 sky130_fd_sc_hd__o211a_1 _12268_ (.A1(_06039_),
    .A2(_05805_),
    .B1(_06044_),
    .C1(_06045_),
    .X(_00381_));
 sky130_fd_sc_hd__nand2_1 _12269_ (.A(_06032_),
    .B(_00974_),
    .Y(_06046_));
 sky130_fd_sc_hd__o211a_1 _12270_ (.A1(_06039_),
    .A2(_05812_),
    .B1(_06044_),
    .C1(_06046_),
    .X(_00382_));
 sky130_fd_sc_hd__nand2_1 _12271_ (.A(_06032_),
    .B(_00999_),
    .Y(_06047_));
 sky130_fd_sc_hd__o211a_1 _12272_ (.A1(_06039_),
    .A2(_05817_),
    .B1(_06044_),
    .C1(_06047_),
    .X(_00383_));
 sky130_fd_sc_hd__nand2_1 _12273_ (.A(_06032_),
    .B(_01024_),
    .Y(_06048_));
 sky130_fd_sc_hd__o211a_1 _12274_ (.A1(_06039_),
    .A2(_05821_),
    .B1(_06044_),
    .C1(_06048_),
    .X(_00384_));
 sky130_fd_sc_hd__nand2_1 _12275_ (.A(_06032_),
    .B(_01049_),
    .Y(_06049_));
 sky130_fd_sc_hd__o211a_1 _12276_ (.A1(_06039_),
    .A2(_05828_),
    .B1(_06044_),
    .C1(_06049_),
    .X(_00385_));
 sky130_fd_sc_hd__nand2_1 _12277_ (.A(_06032_),
    .B(_01075_),
    .Y(_06050_));
 sky130_fd_sc_hd__o211a_1 _12278_ (.A1(_06039_),
    .A2(_05833_),
    .B1(_06044_),
    .C1(_06050_),
    .X(_00386_));
 sky130_fd_sc_hd__nand2_1 _12279_ (.A(_06032_),
    .B(_01101_),
    .Y(_06051_));
 sky130_fd_sc_hd__o211a_1 _12280_ (.A1(_06031_),
    .A2(_05838_),
    .B1(_06044_),
    .C1(_06051_),
    .X(_00387_));
 sky130_fd_sc_hd__and2_1 _12281_ (.A(_02099_),
    .B(_02165_),
    .X(_06052_));
 sky130_fd_sc_hd__and3_1 _12282_ (.A(_00577_),
    .B(_02119_),
    .C(_02120_),
    .X(_06053_));
 sky130_fd_sc_hd__nand2_2 _12283_ (.A(_06052_),
    .B(_06053_),
    .Y(_06054_));
 sky130_fd_sc_hd__buf_2 _12284_ (.A(_06054_),
    .X(_06055_));
 sky130_fd_sc_hd__nand2_1 _12285_ (.A(_06055_),
    .B(_01170_),
    .Y(_06056_));
 sky130_fd_sc_hd__o211a_1 _12286_ (.A1(\R3[0] ),
    .A2(_06055_),
    .B1(_06044_),
    .C1(_06056_),
    .X(_00388_));
 sky130_fd_sc_hd__nand2_1 _12287_ (.A(_06055_),
    .B(_00700_),
    .Y(_06057_));
 sky130_fd_sc_hd__o211a_1 _12288_ (.A1(\R3[1] ),
    .A2(_06055_),
    .B1(_06044_),
    .C1(_06057_),
    .X(_00389_));
 sky130_fd_sc_hd__inv_2 _12289_ (.A(_06054_),
    .Y(_06058_));
 sky130_fd_sc_hd__nand2_1 _12290_ (.A(_06058_),
    .B(\R2[0] ),
    .Y(_06059_));
 sky130_fd_sc_hd__nand2_1 _12291_ (.A(_06055_),
    .B(\result_reg_set[2] ),
    .Y(_06060_));
 sky130_fd_sc_hd__a21oi_1 _12292_ (.A1(_06059_),
    .A2(_06060_),
    .B1(_02116_),
    .Y(_00390_));
 sky130_fd_sc_hd__nand2_1 _12293_ (.A(_06058_),
    .B(\R2[1] ),
    .Y(_06061_));
 sky130_fd_sc_hd__nand2_1 _12294_ (.A(_06055_),
    .B(\result_reg_set[3] ),
    .Y(_06062_));
 sky130_fd_sc_hd__a21oi_1 _12295_ (.A1(_06061_),
    .A2(_06062_),
    .B1(_02116_),
    .Y(_00391_));
 sky130_fd_sc_hd__buf_2 _12296_ (.A(_06058_),
    .X(_06063_));
 sky130_fd_sc_hd__o221a_1 _12297_ (.A1(_05766_),
    .A2(_03172_),
    .B1(_01959_),
    .B2(_02126_),
    .C1(_03175_),
    .X(_06064_));
 sky130_fd_sc_hd__nand2_1 _12298_ (.A(_06063_),
    .B(_06064_),
    .Y(_06065_));
 sky130_fd_sc_hd__o211a_1 _12299_ (.A1(\result_reg_set[4] ),
    .A2(_06063_),
    .B1(_06044_),
    .C1(_06065_),
    .X(_00392_));
 sky130_fd_sc_hd__clkbuf_4 _12300_ (.A(_01148_),
    .X(_06066_));
 sky130_fd_sc_hd__o221a_1 _12301_ (.A1(_05766_),
    .A2(_03131_),
    .B1(_00669_),
    .B2(_02126_),
    .C1(_03144_),
    .X(_06067_));
 sky130_fd_sc_hd__nand2_1 _12302_ (.A(_06063_),
    .B(_06067_),
    .Y(_06068_));
 sky130_fd_sc_hd__o211a_1 _12303_ (.A1(\result_reg_set[5] ),
    .A2(_06063_),
    .B1(_06066_),
    .C1(_06068_),
    .X(_00393_));
 sky130_fd_sc_hd__o221a_1 _12304_ (.A1(_00681_),
    .A2(_02311_),
    .B1(_03094_),
    .B2(_02139_),
    .C1(_03105_),
    .X(_06069_));
 sky130_fd_sc_hd__nand2_1 _12305_ (.A(_06058_),
    .B(_06069_),
    .Y(_06070_));
 sky130_fd_sc_hd__o211a_1 _12306_ (.A1(\result_reg_set[6] ),
    .A2(_06063_),
    .B1(_06066_),
    .C1(_06070_),
    .X(_00394_));
 sky130_fd_sc_hd__o221a_1 _12307_ (.A1(_00671_),
    .A2(_02311_),
    .B1(_01990_),
    .B2(_02139_),
    .C1(_03075_),
    .X(_06071_));
 sky130_fd_sc_hd__nand2_1 _12308_ (.A(_06058_),
    .B(_06071_),
    .Y(_06072_));
 sky130_fd_sc_hd__o211a_1 _12309_ (.A1(\result_reg_set[7] ),
    .A2(_06063_),
    .B1(_06066_),
    .C1(_06072_),
    .X(_00395_));
 sky130_fd_sc_hd__o21ai_1 _12310_ (.A1(_05766_),
    .A2(_01959_),
    .B1(_03834_),
    .Y(_06073_));
 sky130_fd_sc_hd__nand2_1 _12311_ (.A(_06055_),
    .B(_01390_),
    .Y(_06074_));
 sky130_fd_sc_hd__o211a_1 _12312_ (.A1(_06073_),
    .A2(_06055_),
    .B1(_06066_),
    .C1(_06074_),
    .X(_00396_));
 sky130_fd_sc_hd__o21ai_1 _12313_ (.A1(_05766_),
    .A2(_00669_),
    .B1(_03857_),
    .Y(_06075_));
 sky130_fd_sc_hd__nand2_1 _12314_ (.A(_06055_),
    .B(_00930_),
    .Y(_06076_));
 sky130_fd_sc_hd__o211a_1 _12315_ (.A1(_06075_),
    .A2(_06055_),
    .B1(_06066_),
    .C1(_06076_),
    .X(_00397_));
 sky130_fd_sc_hd__nor2_1 _12316_ (.A(_00956_),
    .B(_06058_),
    .Y(_06077_));
 sky130_fd_sc_hd__nor2_1 _12317_ (.A(_05766_),
    .B(_06059_),
    .Y(_06078_));
 sky130_fd_sc_hd__o21a_1 _12318_ (.A1(_06077_),
    .A2(_06078_),
    .B1(_02125_),
    .X(_00398_));
 sky130_fd_sc_hd__nor2_1 _12319_ (.A(_01447_),
    .B(_06058_),
    .Y(_06079_));
 sky130_fd_sc_hd__nor2_1 _12320_ (.A(_05766_),
    .B(_06061_),
    .Y(_06080_));
 sky130_fd_sc_hd__o21a_1 _12321_ (.A1(_06079_),
    .A2(_06080_),
    .B1(_02125_),
    .X(_00399_));
 sky130_fd_sc_hd__a221o_1 _12322_ (.A1(\R3[0] ),
    .A2(_05744_),
    .B1(_00498_),
    .B2(_05745_),
    .C1(_06054_),
    .X(_06081_));
 sky130_fd_sc_hd__o211a_1 _12323_ (.A1(\result_reg_set[12] ),
    .A2(_06063_),
    .B1(_06066_),
    .C1(_06081_),
    .X(_00400_));
 sky130_fd_sc_hd__a221o_1 _12324_ (.A1(\R1[1] ),
    .A2(_05745_),
    .B1(\R3[1] ),
    .B2(_05744_),
    .C1(_06054_),
    .X(_06082_));
 sky130_fd_sc_hd__o211a_1 _12325_ (.A1(\result_reg_set[13] ),
    .A2(_06063_),
    .B1(_06066_),
    .C1(_06082_),
    .X(_00401_));
 sky130_fd_sc_hd__a221o_1 _12326_ (.A1(\R2[0] ),
    .A2(_05744_),
    .B1(\im_reg[6] ),
    .B2(_05745_),
    .C1(_06054_),
    .X(_06083_));
 sky130_fd_sc_hd__o211a_1 _12327_ (.A1(\result_reg_set[14] ),
    .A2(_06063_),
    .B1(_06066_),
    .C1(_06083_),
    .X(_00402_));
 sky130_fd_sc_hd__a221o_1 _12328_ (.A1(\im_reg[7] ),
    .A2(_05745_),
    .B1(\R2[1] ),
    .B2(_05744_),
    .C1(_06054_),
    .X(_06084_));
 sky130_fd_sc_hd__o211a_1 _12329_ (.A1(\result_reg_set[15] ),
    .A2(_06063_),
    .B1(_06066_),
    .C1(_06084_),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_1 _12330_ (.A0(\R3[1] ),
    .A1(net26),
    .S(\current_state[2] ),
    .X(_06085_));
 sky130_fd_sc_hd__and2_1 _12331_ (.A(_06085_),
    .B(_01532_),
    .X(_06086_));
 sky130_fd_sc_hd__clkbuf_1 _12332_ (.A(_06086_),
    .X(_00404_));
 sky130_fd_sc_hd__and2_1 _12333_ (.A(_01529_),
    .B(_01532_),
    .X(_06087_));
 sky130_fd_sc_hd__clkbuf_1 _12334_ (.A(_06087_),
    .X(_00405_));
 sky130_fd_sc_hd__and2_1 _12335_ (.A(_01534_),
    .B(_01532_),
    .X(_06088_));
 sky130_fd_sc_hd__clkbuf_1 _12336_ (.A(_06088_),
    .X(_00406_));
 sky130_fd_sc_hd__mux2_1 _12337_ (.A0(\im_reg[6] ),
    .A1(net31),
    .S(_01146_),
    .X(_06089_));
 sky130_fd_sc_hd__and2_1 _12338_ (.A(_06089_),
    .B(_01532_),
    .X(_06090_));
 sky130_fd_sc_hd__clkbuf_1 _12339_ (.A(_06090_),
    .X(_00407_));
 sky130_fd_sc_hd__mux2_1 _12340_ (.A0(\im_reg[7] ),
    .A1(net32),
    .S(_01146_),
    .X(_06091_));
 sky130_fd_sc_hd__and2_1 _12341_ (.A(_06091_),
    .B(_01532_),
    .X(_06092_));
 sky130_fd_sc_hd__clkbuf_1 _12342_ (.A(_06092_),
    .X(_00408_));
 sky130_fd_sc_hd__mux2_1 _12343_ (.A0(\im_reg[8] ),
    .A1(net33),
    .S(_01146_),
    .X(_06093_));
 sky130_fd_sc_hd__and2_1 _12344_ (.A(_06093_),
    .B(_01532_),
    .X(_06094_));
 sky130_fd_sc_hd__clkbuf_1 _12345_ (.A(_06094_),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_1 _12346_ (.A0(\im_reg[9] ),
    .A1(net34),
    .S(_01146_),
    .X(_06095_));
 sky130_fd_sc_hd__and2_1 _12347_ (.A(_06095_),
    .B(_01532_),
    .X(_06096_));
 sky130_fd_sc_hd__clkbuf_1 _12348_ (.A(_06096_),
    .X(_00410_));
 sky130_fd_sc_hd__buf_2 _12349_ (.A(_01146_),
    .X(_06097_));
 sky130_fd_sc_hd__nor2_1 _12350_ (.A(net24),
    .B(net25),
    .Y(_06098_));
 sky130_fd_sc_hd__nand2_1 _12351_ (.A(net22),
    .B(net21),
    .Y(_06099_));
 sky130_fd_sc_hd__inv_2 _12352_ (.A(net23),
    .Y(_06100_));
 sky130_fd_sc_hd__a31o_1 _12353_ (.A1(_06098_),
    .A2(_06099_),
    .A3(_06100_),
    .B1(_06267_),
    .X(_06101_));
 sky130_fd_sc_hd__o211a_1 _12354_ (.A1(_06097_),
    .A2(CMD_addition),
    .B1(_06066_),
    .C1(_06101_),
    .X(_00411_));
 sky130_fd_sc_hd__clkbuf_4 _12355_ (.A(_01146_),
    .X(_06102_));
 sky130_fd_sc_hd__nor2_1 _12356_ (.A(_06102_),
    .B(_00528_),
    .Y(_06103_));
 sky130_fd_sc_hd__nand2_1 _12357_ (.A(net22),
    .B(net23),
    .Y(_06104_));
 sky130_fd_sc_hd__inv_2 _12358_ (.A(_06104_),
    .Y(_06105_));
 sky130_fd_sc_hd__inv_2 _12359_ (.A(_06098_),
    .Y(_06106_));
 sky130_fd_sc_hd__nor2_1 _12360_ (.A(net22),
    .B(net21),
    .Y(_06107_));
 sky130_fd_sc_hd__a31o_1 _12361_ (.A1(_06107_),
    .A2(_06100_),
    .A3(_06253_),
    .B1(_06098_),
    .X(_06108_));
 sky130_fd_sc_hd__o211a_1 _12362_ (.A1(_06105_),
    .A2(_06106_),
    .B1(_06102_),
    .C1(_06108_),
    .X(_06109_));
 sky130_fd_sc_hd__o21a_1 _12363_ (.A1(_06103_),
    .A2(_06109_),
    .B1(_02125_),
    .X(_00412_));
 sky130_fd_sc_hd__a211o_1 _12364_ (.A1(_06100_),
    .A2(_06099_),
    .B1(_06105_),
    .C1(_06106_),
    .X(_06110_));
 sky130_fd_sc_hd__nand2_1 _12365_ (.A(_06110_),
    .B(_06097_),
    .Y(_06111_));
 sky130_fd_sc_hd__o211a_1 _12366_ (.A1(_06097_),
    .A2(_02160_),
    .B1(_04827_),
    .C1(_06111_),
    .X(_00413_));
 sky130_fd_sc_hd__nor2_2 _12367_ (.A(net22),
    .B(net23),
    .Y(_06112_));
 sky130_fd_sc_hd__inv_2 _12368_ (.A(_06112_),
    .Y(_06113_));
 sky130_fd_sc_hd__inv_2 _12369_ (.A(net22),
    .Y(_06114_));
 sky130_fd_sc_hd__nor2_1 _12370_ (.A(net23),
    .B(_06114_),
    .Y(_06115_));
 sky130_fd_sc_hd__nor2_2 _12371_ (.A(net20),
    .B(net21),
    .Y(_06116_));
 sky130_fd_sc_hd__nand2_2 _12372_ (.A(_06115_),
    .B(_06116_),
    .Y(_06117_));
 sky130_fd_sc_hd__a311o_1 _12373_ (.A1(net24),
    .A2(_06113_),
    .A3(_06117_),
    .B1(net25),
    .C1(_06108_),
    .X(_06118_));
 sky130_fd_sc_hd__nor2_1 _12374_ (.A(_06102_),
    .B(_04830_),
    .Y(_06119_));
 sky130_fd_sc_hd__a211oi_2 _12375_ (.A1(_06118_),
    .A2(_06102_),
    .B1(_02115_),
    .C1(_06119_),
    .Y(_00414_));
 sky130_fd_sc_hd__or4_1 _12376_ (.A(net22),
    .B(net25),
    .C(_06254_),
    .D(_06256_),
    .X(_06120_));
 sky130_fd_sc_hd__nand2_1 _12377_ (.A(_06120_),
    .B(_06097_),
    .Y(_06121_));
 sky130_fd_sc_hd__o211a_1 _12378_ (.A1(_06097_),
    .A2(CMD_logic_shift_right),
    .B1(_04827_),
    .C1(_06121_),
    .X(_00415_));
 sky130_fd_sc_hd__inv_2 _12379_ (.A(net24),
    .Y(_06122_));
 sky130_fd_sc_hd__nor2_2 _12380_ (.A(net25),
    .B(_06122_),
    .Y(_06123_));
 sky130_fd_sc_hd__nand2_2 _12381_ (.A(_06123_),
    .B(\current_state[2] ),
    .Y(_06124_));
 sky130_fd_sc_hd__or4_1 _12382_ (.A(_06114_),
    .B(net23),
    .C(_06116_),
    .D(_06124_),
    .X(_06125_));
 sky130_fd_sc_hd__buf_2 _12383_ (.A(_06267_),
    .X(_06126_));
 sky130_fd_sc_hd__nand2_1 _12384_ (.A(_06126_),
    .B(_02118_),
    .Y(_06127_));
 sky130_fd_sc_hd__a21oi_1 _12385_ (.A1(_06125_),
    .A2(_06127_),
    .B1(_02116_),
    .Y(_00416_));
 sky130_fd_sc_hd__nor2_2 _12386_ (.A(net22),
    .B(_06100_),
    .Y(_06128_));
 sky130_fd_sc_hd__nand2_1 _12387_ (.A(_06128_),
    .B(_06256_),
    .Y(_06129_));
 sky130_fd_sc_hd__inv_2 _12388_ (.A(_06123_),
    .Y(_06130_));
 sky130_fd_sc_hd__inv_2 _12389_ (.A(net20),
    .Y(_06131_));
 sky130_fd_sc_hd__and2_1 _12390_ (.A(_06131_),
    .B(net21),
    .X(_06132_));
 sky130_fd_sc_hd__nand2_1 _12391_ (.A(_06132_),
    .B(_06105_),
    .Y(_06133_));
 sky130_fd_sc_hd__nor2_1 _12392_ (.A(_06130_),
    .B(_06133_),
    .Y(_06134_));
 sky130_fd_sc_hd__o21bai_1 _12393_ (.A1(_06254_),
    .A2(_06257_),
    .B1_N(_06134_),
    .Y(_06135_));
 sky130_fd_sc_hd__a2111oi_1 _12394_ (.A1(_06104_),
    .A2(_06129_),
    .B1(_06122_),
    .C1(net25),
    .D1(_06135_),
    .Y(_06136_));
 sky130_fd_sc_hd__nand2_1 _12395_ (.A(_06126_),
    .B(_00547_),
    .Y(_06137_));
 sky130_fd_sc_hd__o211a_1 _12396_ (.A1(_06126_),
    .A2(_06136_),
    .B1(_04827_),
    .C1(_06137_),
    .X(_00417_));
 sky130_fd_sc_hd__nor2_1 _12397_ (.A(net24),
    .B(_06253_),
    .Y(_06138_));
 sky130_fd_sc_hd__inv_2 _12398_ (.A(_06138_),
    .Y(_06139_));
 sky130_fd_sc_hd__inv_2 _12399_ (.A(_06116_),
    .Y(_06140_));
 sky130_fd_sc_hd__nor2_1 _12400_ (.A(_06113_),
    .B(_06140_),
    .Y(_06141_));
 sky130_fd_sc_hd__inv_2 _12401_ (.A(_06141_),
    .Y(_06142_));
 sky130_fd_sc_hd__nor2_1 _12402_ (.A(_06139_),
    .B(_06142_),
    .Y(_06143_));
 sky130_fd_sc_hd__a211o_1 _12403_ (.A1(_06135_),
    .A2(_06253_),
    .B1(_06267_),
    .C1(_06143_),
    .X(_06144_));
 sky130_fd_sc_hd__o211a_1 _12404_ (.A1(_06097_),
    .A2(_00545_),
    .B1(_04827_),
    .C1(_06144_),
    .X(_00418_));
 sky130_fd_sc_hd__nor2_1 _12405_ (.A(_06102_),
    .B(_00578_),
    .Y(_06145_));
 sky130_fd_sc_hd__and4_1 _12406_ (.A(_06140_),
    .B(_06138_),
    .C(_06112_),
    .D(_01146_),
    .X(_06146_));
 sky130_fd_sc_hd__o21a_1 _12407_ (.A1(_06145_),
    .A2(_06146_),
    .B1(_02125_),
    .X(_00419_));
 sky130_fd_sc_hd__nand2_1 _12408_ (.A(_06132_),
    .B(_06115_),
    .Y(_06147_));
 sky130_fd_sc_hd__a41o_1 _12409_ (.A1(_06147_),
    .A2(_06257_),
    .A3(_06100_),
    .A4(_06122_),
    .B1(_06253_),
    .X(_06148_));
 sky130_fd_sc_hd__nand2_2 _12410_ (.A(_06128_),
    .B(_06116_),
    .Y(_06149_));
 sky130_fd_sc_hd__a21o_1 _12411_ (.A1(_06149_),
    .A2(net23),
    .B1(_06139_),
    .X(_06150_));
 sky130_fd_sc_hd__nand2_1 _12412_ (.A(_06150_),
    .B(net25),
    .Y(_06151_));
 sky130_fd_sc_hd__or3b_1 _12413_ (.A(_06266_),
    .B(_06148_),
    .C_N(_06151_),
    .X(_06152_));
 sky130_fd_sc_hd__nand2_1 _12414_ (.A(_06126_),
    .B(CMD_load),
    .Y(_06153_));
 sky130_fd_sc_hd__a21oi_1 _12415_ (.A1(_06152_),
    .A2(_06153_),
    .B1(_02116_),
    .Y(_00420_));
 sky130_fd_sc_hd__a21oi_1 _12416_ (.A1(_06104_),
    .A2(_06122_),
    .B1(_06253_),
    .Y(_06154_));
 sky130_fd_sc_hd__or3_1 _12417_ (.A(_06266_),
    .B(_06154_),
    .C(_06151_),
    .X(_06155_));
 sky130_fd_sc_hd__nand2_1 _12418_ (.A(_06126_),
    .B(CMD_store),
    .Y(_06156_));
 sky130_fd_sc_hd__a21oi_1 _12419_ (.A1(_06155_),
    .A2(_06156_),
    .B1(_02116_),
    .Y(_00421_));
 sky130_fd_sc_hd__nand2_1 _12420_ (.A(_06256_),
    .B(_06105_),
    .Y(_06157_));
 sky130_fd_sc_hd__and3_1 _12421_ (.A(_06154_),
    .B(_06122_),
    .C(_06157_),
    .X(_06158_));
 sky130_fd_sc_hd__nand2_1 _12422_ (.A(_06126_),
    .B(_00576_),
    .Y(_06159_));
 sky130_fd_sc_hd__o211a_1 _12423_ (.A1(_06126_),
    .A2(_06158_),
    .B1(_04827_),
    .C1(_06159_),
    .X(_00422_));
 sky130_fd_sc_hd__or3_1 _12424_ (.A(net24),
    .B(_06266_),
    .C(_06253_),
    .X(_06160_));
 sky130_fd_sc_hd__or2_1 _12425_ (.A(_06117_),
    .B(_06160_),
    .X(_06161_));
 sky130_fd_sc_hd__nand2_1 _12426_ (.A(_06126_),
    .B(CMD_loopjump),
    .Y(_06162_));
 sky130_fd_sc_hd__a21oi_1 _12427_ (.A1(_06161_),
    .A2(_06162_),
    .B1(_02116_),
    .Y(_00423_));
 sky130_fd_sc_hd__nor2_1 _12428_ (.A(_06102_),
    .B(_01962_),
    .Y(_06163_));
 sky130_fd_sc_hd__nor2_1 _12429_ (.A(net21),
    .B(_06131_),
    .Y(_06164_));
 sky130_fd_sc_hd__nand2_1 _12430_ (.A(_06115_),
    .B(_06164_),
    .Y(_06165_));
 sky130_fd_sc_hd__nor2_1 _12431_ (.A(_06165_),
    .B(_06160_),
    .Y(_06166_));
 sky130_fd_sc_hd__o21a_1 _12432_ (.A1(_06163_),
    .A2(_06166_),
    .B1(_02125_),
    .X(_00424_));
 sky130_fd_sc_hd__nand2_1 _12433_ (.A(_06164_),
    .B(_06112_),
    .Y(_06167_));
 sky130_fd_sc_hd__a21o_1 _12434_ (.A1(_06165_),
    .A2(_06149_),
    .B1(_06124_),
    .X(_06168_));
 sky130_fd_sc_hd__o221a_1 _12435_ (.A1(_01146_),
    .A2(_01554_),
    .B1(_06167_),
    .B2(_06160_),
    .C1(_06168_),
    .X(_06169_));
 sky130_fd_sc_hd__nor2_1 _12436_ (.A(_06255_),
    .B(_06113_),
    .Y(_06170_));
 sky130_fd_sc_hd__inv_2 _12437_ (.A(_06170_),
    .Y(_06171_));
 sky130_fd_sc_hd__nand2_1 _12438_ (.A(_06164_),
    .B(_06128_),
    .Y(_06172_));
 sky130_fd_sc_hd__a31o_1 _12439_ (.A1(_06171_),
    .A2(_06157_),
    .A3(_06172_),
    .B1(_06106_),
    .X(_06173_));
 sky130_fd_sc_hd__nor2_1 _12440_ (.A(_06104_),
    .B(_06140_),
    .Y(_06174_));
 sky130_fd_sc_hd__nand2_1 _12441_ (.A(_06147_),
    .B(_06172_),
    .Y(_06175_));
 sky130_fd_sc_hd__o21ai_1 _12442_ (.A1(_06174_),
    .A2(_06175_),
    .B1(_06138_),
    .Y(_06176_));
 sky130_fd_sc_hd__a21o_1 _12443_ (.A1(_06173_),
    .A2(_06176_),
    .B1(_06267_),
    .X(_06177_));
 sky130_fd_sc_hd__a21oi_1 _12444_ (.A1(_06169_),
    .A2(_06177_),
    .B1(_02116_),
    .Y(_00425_));
 sky130_fd_sc_hd__inv_2 _12445_ (.A(_06174_),
    .Y(_06178_));
 sky130_fd_sc_hd__a31oi_1 _12446_ (.A1(_06142_),
    .A2(_06178_),
    .A3(_06147_),
    .B1(_06106_),
    .Y(_06179_));
 sky130_fd_sc_hd__a311o_1 _12447_ (.A1(_06123_),
    .A2(_06128_),
    .A3(_06256_),
    .B1(_06267_),
    .C1(_06134_),
    .X(_06180_));
 sky130_fd_sc_hd__o221a_1 _12448_ (.A1(_06097_),
    .A2(_05904_),
    .B1(_06179_),
    .B2(_06180_),
    .C1(_02101_),
    .X(_00426_));
 sky130_fd_sc_hd__nand2_1 _12449_ (.A(_06132_),
    .B(_06112_),
    .Y(_06181_));
 sky130_fd_sc_hd__nor2_1 _12450_ (.A(_06130_),
    .B(_06181_),
    .Y(_06182_));
 sky130_fd_sc_hd__nand2_1 _12451_ (.A(_06126_),
    .B(_00626_),
    .Y(_06183_));
 sky130_fd_sc_hd__o211a_1 _12452_ (.A1(_06126_),
    .A2(_06182_),
    .B1(_04827_),
    .C1(_06183_),
    .X(_00427_));
 sky130_fd_sc_hd__nand2_1 _12453_ (.A(_06267_),
    .B(Him),
    .Y(_06184_));
 sky130_fd_sc_hd__a21oi_1 _12454_ (.A1(_06177_),
    .A2(_06184_),
    .B1(_02650_),
    .Y(_00428_));
 sky130_fd_sc_hd__a2bb2o_1 _12455_ (.A1_N(_06139_),
    .A2_N(_06181_),
    .B1(_06123_),
    .B2(_06175_),
    .X(_06185_));
 sky130_fd_sc_hd__nand2_1 _12456_ (.A(_06132_),
    .B(_06128_),
    .Y(_06186_));
 sky130_fd_sc_hd__nand2_1 _12457_ (.A(_06186_),
    .B(_06117_),
    .Y(_06187_));
 sky130_fd_sc_hd__nand2_1 _12458_ (.A(_06164_),
    .B(_06105_),
    .Y(_06188_));
 sky130_fd_sc_hd__inv_2 _12459_ (.A(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__nor2_1 _12460_ (.A(net23),
    .B(_06257_),
    .Y(_06190_));
 sky130_fd_sc_hd__nor2_1 _12461_ (.A(_06189_),
    .B(_06190_),
    .Y(_06191_));
 sky130_fd_sc_hd__nand2_1 _12462_ (.A(_06191_),
    .B(_06186_),
    .Y(_06192_));
 sky130_fd_sc_hd__a31o_1 _12463_ (.A1(_06123_),
    .A2(_06112_),
    .A3(_06116_),
    .B1(_06266_),
    .X(_06193_));
 sky130_fd_sc_hd__a221o_1 _12464_ (.A1(_06098_),
    .A2(_06187_),
    .B1(_06192_),
    .B2(_06138_),
    .C1(_06193_),
    .X(_06194_));
 sky130_fd_sc_hd__o221a_1 _12465_ (.A1(_06097_),
    .A2(_00585_),
    .B1(_06185_),
    .B2(_06194_),
    .C1(_02101_),
    .X(_00429_));
 sky130_fd_sc_hd__a21oi_1 _12466_ (.A1(_06191_),
    .A2(_06167_),
    .B1(_06106_),
    .Y(_06195_));
 sky130_fd_sc_hd__nand2_1 _12467_ (.A(_06178_),
    .B(_06157_),
    .Y(_06196_));
 sky130_fd_sc_hd__a21o_1 _12468_ (.A1(_06196_),
    .A2(_06123_),
    .B1(_06267_),
    .X(_06197_));
 sky130_fd_sc_hd__o221a_1 _12469_ (.A1(_06097_),
    .A2(Oreg2),
    .B1(_06195_),
    .B2(_06197_),
    .C1(_02101_),
    .X(_00430_));
 sky130_fd_sc_hd__o22a_1 _12470_ (.A1(_06102_),
    .A2(_00647_),
    .B1(_06124_),
    .B2(_06171_),
    .X(_06198_));
 sky130_fd_sc_hd__nor2_1 _12471_ (.A(_02116_),
    .B(_06198_),
    .Y(_00431_));
 sky130_fd_sc_hd__o211a_1 _12472_ (.A1(_06097_),
    .A2(Oim),
    .B1(_04827_),
    .C1(_06194_),
    .X(_00432_));
 sky130_fd_sc_hd__a31o_1 _12473_ (.A1(_06133_),
    .A2(_06149_),
    .A3(_06129_),
    .B1(_06139_),
    .X(_06199_));
 sky130_fd_sc_hd__and2_1 _12474_ (.A(_06165_),
    .B(_06129_),
    .X(_06200_));
 sky130_fd_sc_hd__o22a_1 _12475_ (.A1(_06130_),
    .A2(_06167_),
    .B1(_06106_),
    .B2(_06200_),
    .X(_06201_));
 sky130_fd_sc_hd__and3_1 _12476_ (.A(_06199_),
    .B(_01146_),
    .C(_06201_),
    .X(_06202_));
 sky130_fd_sc_hd__nand2_1 _12477_ (.A(_06190_),
    .B(_06123_),
    .Y(_06203_));
 sky130_fd_sc_hd__o221a_1 _12478_ (.A1(_06130_),
    .A2(_06186_),
    .B1(_06139_),
    .B2(_06171_),
    .C1(_06203_),
    .X(_06204_));
 sky130_fd_sc_hd__a221o_1 _12479_ (.A1(_06267_),
    .A2(_00582_),
    .B1(_06202_),
    .B2(_06204_),
    .C1(_05775_),
    .X(_06205_));
 sky130_fd_sc_hd__inv_2 _12480_ (.A(_06205_),
    .Y(_00433_));
 sky130_fd_sc_hd__a31oi_1 _12481_ (.A1(_06181_),
    .A2(_06133_),
    .A3(_06149_),
    .B1(_06106_),
    .Y(_06206_));
 sky130_fd_sc_hd__a211o_1 _12482_ (.A1(_06123_),
    .A2(_06189_),
    .B1(_06267_),
    .C1(_06143_),
    .X(_06207_));
 sky130_fd_sc_hd__o221a_1 _12483_ (.A1(_06102_),
    .A2(Qreg2),
    .B1(_06206_),
    .B2(_06207_),
    .C1(_02101_),
    .X(_00434_));
 sky130_fd_sc_hd__o22a_1 _12484_ (.A1(_06102_),
    .A2(_00620_),
    .B1(_06117_),
    .B2(_06124_),
    .X(_06208_));
 sky130_fd_sc_hd__nor2_1 _12485_ (.A(_02116_),
    .B(_06208_),
    .Y(_00435_));
 sky130_fd_sc_hd__o21ai_1 _12486_ (.A1(_06102_),
    .A2(Qim),
    .B1(_04827_),
    .Y(_06209_));
 sky130_fd_sc_hd__nor2_1 _12487_ (.A(_06209_),
    .B(_06202_),
    .Y(_00436_));
 sky130_fd_sc_hd__and2_1 _12488_ (.A(_01147_),
    .B(_05134_),
    .X(_06210_));
 sky130_fd_sc_hd__clkbuf_1 _12489_ (.A(_06210_),
    .X(_00437_));
 sky130_fd_sc_hd__and2_1 _12490_ (.A(_01151_),
    .B(_05134_),
    .X(_06211_));
 sky130_fd_sc_hd__clkbuf_1 _12491_ (.A(_06211_),
    .X(_00438_));
 sky130_fd_sc_hd__and2_1 _12492_ (.A(_01531_),
    .B(_05134_),
    .X(_06212_));
 sky130_fd_sc_hd__clkbuf_1 _12493_ (.A(_06212_),
    .X(_00439_));
 sky130_fd_sc_hd__and2_1 _12494_ (.A(_01527_),
    .B(_05134_),
    .X(_06213_));
 sky130_fd_sc_hd__clkbuf_1 _12495_ (.A(_06213_),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _12496_ (.A0(\R3[0] ),
    .A1(net17),
    .S(\current_state[2] ),
    .X(_06214_));
 sky130_fd_sc_hd__and2_1 _12497_ (.A(_06214_),
    .B(_01532_),
    .X(_06215_));
 sky130_fd_sc_hd__clkbuf_1 _12498_ (.A(_06215_),
    .X(_00441_));
 sky130_fd_sc_hd__and4b_1 _12499_ (.A_N(\current_state[1] ),
    .B(_06271_),
    .C(_06269_),
    .D(_00631_),
    .X(_06216_));
 sky130_fd_sc_hd__and3_1 _12500_ (.A(_06216_),
    .B(_06266_),
    .C(_06263_),
    .X(_06217_));
 sky130_fd_sc_hd__nand2_4 _12501_ (.A(_06217_),
    .B(_06258_),
    .Y(_06218_));
 sky130_fd_sc_hd__inv_2 _12502_ (.A(_06218_),
    .Y(_06219_));
 sky130_fd_sc_hd__clkbuf_4 _12503_ (.A(_06219_),
    .X(_06220_));
 sky130_fd_sc_hd__clkbuf_4 _12504_ (.A(_06259_),
    .X(_06221_));
 sky130_fd_sc_hd__or2_1 _12505_ (.A(\next_PC[0] ),
    .B(_06218_),
    .X(_06222_));
 sky130_fd_sc_hd__o211a_1 _12506_ (.A1(net65),
    .A2(_06220_),
    .B1(_06221_),
    .C1(_06222_),
    .X(_00442_));
 sky130_fd_sc_hd__or2_1 _12507_ (.A(\next_PC[1] ),
    .B(_06218_),
    .X(_06223_));
 sky130_fd_sc_hd__o211a_1 _12508_ (.A1(net66),
    .A2(_06220_),
    .B1(_06221_),
    .C1(_06223_),
    .X(_00443_));
 sky130_fd_sc_hd__or2_1 _12509_ (.A(\next_PC[2] ),
    .B(_06218_),
    .X(_06224_));
 sky130_fd_sc_hd__o211a_1 _12510_ (.A1(net67),
    .A2(_06220_),
    .B1(_06221_),
    .C1(_06224_),
    .X(_00444_));
 sky130_fd_sc_hd__nand2_1 _12511_ (.A(_06219_),
    .B(_00490_),
    .Y(_06225_));
 sky130_fd_sc_hd__o211a_1 _12512_ (.A1(net68),
    .A2(_06220_),
    .B1(_06221_),
    .C1(_06225_),
    .X(_00445_));
 sky130_fd_sc_hd__or2_1 _12513_ (.A(\next_PC[4] ),
    .B(_06218_),
    .X(_06226_));
 sky130_fd_sc_hd__o211a_1 _12514_ (.A1(net69),
    .A2(_06220_),
    .B1(_06221_),
    .C1(_06226_),
    .X(_00446_));
 sky130_fd_sc_hd__nand2_1 _12515_ (.A(_06219_),
    .B(_00500_),
    .Y(_06227_));
 sky130_fd_sc_hd__o211a_1 _12516_ (.A1(net70),
    .A2(_06220_),
    .B1(_06221_),
    .C1(_06227_),
    .X(_00447_));
 sky130_fd_sc_hd__nand2_1 _12517_ (.A(_06219_),
    .B(_00506_),
    .Y(_06228_));
 sky130_fd_sc_hd__o211a_1 _12518_ (.A1(net71),
    .A2(_06220_),
    .B1(_06221_),
    .C1(_06228_),
    .X(_00448_));
 sky130_fd_sc_hd__or2_1 _12519_ (.A(\next_PC[7] ),
    .B(_06218_),
    .X(_06229_));
 sky130_fd_sc_hd__o211a_1 _12520_ (.A1(net72),
    .A2(_06220_),
    .B1(_06221_),
    .C1(_06229_),
    .X(_00449_));
 sky130_fd_sc_hd__nand2_1 _12521_ (.A(_06219_),
    .B(_00515_),
    .Y(_06230_));
 sky130_fd_sc_hd__o211a_1 _12522_ (.A1(net73),
    .A2(_06220_),
    .B1(_06221_),
    .C1(_06230_),
    .X(_00450_));
 sky130_fd_sc_hd__or2_1 _12523_ (.A(\next_PC[9] ),
    .B(_06218_),
    .X(_06231_));
 sky130_fd_sc_hd__o211a_1 _12524_ (.A1(net74),
    .A2(_06220_),
    .B1(_06221_),
    .C1(_06231_),
    .X(_00451_));
 sky130_fd_sc_hd__or2_1 _12525_ (.A(_00685_),
    .B(_01126_),
    .X(_06232_));
 sky130_fd_sc_hd__clkbuf_4 _12526_ (.A(_06232_),
    .X(_06233_));
 sky130_fd_sc_hd__clkbuf_8 _12527_ (.A(_06233_),
    .X(_06234_));
 sky130_fd_sc_hd__mux2_1 _12528_ (.A0(_00668_),
    .A1(\Qset[3][0] ),
    .S(_06234_),
    .X(_06235_));
 sky130_fd_sc_hd__clkbuf_1 _12529_ (.A(_06235_),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _12530_ (.A0(_00722_),
    .A1(\Qset[3][1] ),
    .S(_06234_),
    .X(_06236_));
 sky130_fd_sc_hd__clkbuf_1 _12531_ (.A(_06236_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _12532_ (.A0(_00759_),
    .A1(\Qset[3][2] ),
    .S(_06234_),
    .X(_06237_));
 sky130_fd_sc_hd__clkbuf_1 _12533_ (.A(_06237_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _12534_ (.A0(_00783_),
    .A1(\Qset[3][3] ),
    .S(_06234_),
    .X(_06238_));
 sky130_fd_sc_hd__clkbuf_1 _12535_ (.A(_06238_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _12536_ (.A0(_00809_),
    .A1(\Qset[3][4] ),
    .S(_06234_),
    .X(_06239_));
 sky130_fd_sc_hd__clkbuf_1 _12537_ (.A(_06239_),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _12538_ (.A0(_00854_),
    .A1(\Qset[3][5] ),
    .S(_06234_),
    .X(_06240_));
 sky130_fd_sc_hd__clkbuf_1 _12539_ (.A(_06240_),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _12540_ (.A0(_00878_),
    .A1(\Qset[3][6] ),
    .S(_06234_),
    .X(_06241_));
 sky130_fd_sc_hd__clkbuf_1 _12541_ (.A(_06241_),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_1 _12542_ (.A0(_00904_),
    .A1(\Qset[3][7] ),
    .S(_06234_),
    .X(_06242_));
 sky130_fd_sc_hd__clkbuf_1 _12543_ (.A(_06242_),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _12544_ (.A0(_00927_),
    .A1(\Qset[3][8] ),
    .S(_06234_),
    .X(_06243_));
 sky130_fd_sc_hd__clkbuf_1 _12545_ (.A(_06243_),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _12546_ (.A0(_00953_),
    .A1(\Qset[3][9] ),
    .S(_06234_),
    .X(_06244_));
 sky130_fd_sc_hd__clkbuf_1 _12547_ (.A(_06244_),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _12548_ (.A0(_00979_),
    .A1(\Qset[3][10] ),
    .S(_06233_),
    .X(_06245_));
 sky130_fd_sc_hd__clkbuf_1 _12549_ (.A(_06245_),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _12550_ (.A0(_01004_),
    .A1(\Qset[3][11] ),
    .S(_06233_),
    .X(_06246_));
 sky130_fd_sc_hd__clkbuf_1 _12551_ (.A(_06246_),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _12552_ (.A0(_01029_),
    .A1(\Qset[3][12] ),
    .S(_06233_),
    .X(_06247_));
 sky130_fd_sc_hd__clkbuf_1 _12553_ (.A(_06247_),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _12554_ (.A0(_01054_),
    .A1(\Qset[3][13] ),
    .S(_06233_),
    .X(_06248_));
 sky130_fd_sc_hd__clkbuf_1 _12555_ (.A(_06248_),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _12556_ (.A0(_01080_),
    .A1(\Qset[3][14] ),
    .S(_06233_),
    .X(_06249_));
 sky130_fd_sc_hd__clkbuf_1 _12557_ (.A(_06249_),
    .X(_00466_));
 sky130_fd_sc_hd__mux2_1 _12558_ (.A0(_01106_),
    .A1(\Qset[3][15] ),
    .S(_06233_),
    .X(_06250_));
 sky130_fd_sc_hd__clkbuf_1 _12559_ (.A(_06250_),
    .X(_00467_));
 sky130_fd_sc_hd__and2_1 _12560_ (.A(_06214_),
    .B(_05134_),
    .X(_06251_));
 sky130_fd_sc_hd__clkbuf_1 _12561_ (.A(_06251_),
    .X(_00468_));
 sky130_fd_sc_hd__and2_1 _12562_ (.A(_06085_),
    .B(_05134_),
    .X(_06252_));
 sky130_fd_sc_hd__clkbuf_1 _12563_ (.A(_06252_),
    .X(_00469_));
 sky130_fd_sc_hd__dfxtp_1 _12564_ (.CLK(clknet_leaf_39_clk),
    .D(_00014_),
    .Q(\next_PC[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12565_ (.CLK(clknet_leaf_39_clk),
    .D(_00015_),
    .Q(\next_PC[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12566_ (.CLK(clknet_leaf_38_clk),
    .D(_00016_),
    .Q(\next_PC[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12567_ (.CLK(clknet_leaf_38_clk),
    .D(_00017_),
    .Q(\next_PC[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12568_ (.CLK(clknet_leaf_38_clk),
    .D(_00018_),
    .Q(\next_PC[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12569_ (.CLK(clknet_leaf_38_clk),
    .D(_00019_),
    .Q(\next_PC[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12570_ (.CLK(clknet_leaf_36_clk),
    .D(_00020_),
    .Q(\next_PC[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12571_ (.CLK(clknet_leaf_34_clk),
    .D(_00021_),
    .Q(\next_PC[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12572_ (.CLK(clknet_leaf_34_clk),
    .D(_00022_),
    .Q(\next_PC[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12573_ (.CLK(clknet_leaf_28_clk),
    .D(_00023_),
    .Q(\next_PC[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12574_ (.CLK(clknet_leaf_49_clk),
    .D(_00024_),
    .Q(\Qset[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12575_ (.CLK(clknet_leaf_46_clk),
    .D(_00025_),
    .Q(\Qset[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12576_ (.CLK(clknet_leaf_45_clk),
    .D(_00026_),
    .Q(\Qset[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12577_ (.CLK(clknet_leaf_48_clk),
    .D(_00027_),
    .Q(\Qset[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12578_ (.CLK(clknet_leaf_48_clk),
    .D(_00028_),
    .Q(\Qset[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12579_ (.CLK(clknet_leaf_45_clk),
    .D(_00029_),
    .Q(\Qset[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12580_ (.CLK(clknet_leaf_44_clk),
    .D(_00030_),
    .Q(\Qset[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12581_ (.CLK(clknet_leaf_43_clk),
    .D(_00031_),
    .Q(\Qset[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12582_ (.CLK(clknet_leaf_40_clk),
    .D(_00032_),
    .Q(\Qset[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12583_ (.CLK(clknet_leaf_40_clk),
    .D(_00033_),
    .Q(\Qset[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12584_ (.CLK(clknet_leaf_33_clk),
    .D(_00034_),
    .Q(\Qset[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12585_ (.CLK(clknet_leaf_35_clk),
    .D(_00035_),
    .Q(\Qset[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12586_ (.CLK(clknet_leaf_29_clk),
    .D(_00036_),
    .Q(\Qset[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12587_ (.CLK(clknet_leaf_28_clk),
    .D(_00037_),
    .Q(\Qset[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12588_ (.CLK(clknet_leaf_27_clk),
    .D(_00038_),
    .Q(\Qset[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12589_ (.CLK(clknet_leaf_26_clk),
    .D(_00039_),
    .Q(\Qset[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12590_ (.CLK(clknet_leaf_49_clk),
    .D(_00040_),
    .Q(\Qset[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12591_ (.CLK(clknet_leaf_46_clk),
    .D(_00041_),
    .Q(\Qset[1][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12592_ (.CLK(clknet_leaf_46_clk),
    .D(_00042_),
    .Q(\Qset[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12593_ (.CLK(clknet_leaf_48_clk),
    .D(_00043_),
    .Q(\Qset[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12594_ (.CLK(clknet_leaf_48_clk),
    .D(_00044_),
    .Q(\Qset[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12595_ (.CLK(clknet_leaf_45_clk),
    .D(_00045_),
    .Q(\Qset[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12596_ (.CLK(clknet_leaf_43_clk),
    .D(_00046_),
    .Q(\Qset[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12597_ (.CLK(clknet_leaf_43_clk),
    .D(_00047_),
    .Q(\Qset[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12598_ (.CLK(clknet_leaf_40_clk),
    .D(_00048_),
    .Q(\Qset[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12599_ (.CLK(clknet_leaf_39_clk),
    .D(_00049_),
    .Q(\Qset[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12600_ (.CLK(clknet_leaf_34_clk),
    .D(_00050_),
    .Q(\Qset[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12601_ (.CLK(clknet_leaf_35_clk),
    .D(_00051_),
    .Q(\Qset[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12602_ (.CLK(clknet_leaf_34_clk),
    .D(_00052_),
    .Q(\Qset[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12603_ (.CLK(clknet_leaf_28_clk),
    .D(_00053_),
    .Q(\Qset[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12604_ (.CLK(clknet_leaf_25_clk),
    .D(_00054_),
    .Q(\Qset[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12605_ (.CLK(clknet_leaf_25_clk),
    .D(_00055_),
    .Q(\Qset[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12606_ (.CLK(clknet_leaf_49_clk),
    .D(_00056_),
    .Q(\Qset[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12607_ (.CLK(clknet_leaf_46_clk),
    .D(_00057_),
    .Q(\Qset[2][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12608_ (.CLK(clknet_leaf_46_clk),
    .D(_00058_),
    .Q(\Qset[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12609_ (.CLK(clknet_leaf_48_clk),
    .D(_00059_),
    .Q(\Qset[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12610_ (.CLK(clknet_leaf_48_clk),
    .D(_00060_),
    .Q(\Qset[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12611_ (.CLK(clknet_leaf_45_clk),
    .D(_00061_),
    .Q(\Qset[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12612_ (.CLK(clknet_leaf_43_clk),
    .D(_00062_),
    .Q(\Qset[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12613_ (.CLK(clknet_leaf_43_clk),
    .D(_00063_),
    .Q(\Qset[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12614_ (.CLK(clknet_leaf_40_clk),
    .D(_00064_),
    .Q(\Qset[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12615_ (.CLK(clknet_leaf_39_clk),
    .D(_00065_),
    .Q(\Qset[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12616_ (.CLK(clknet_leaf_35_clk),
    .D(_00066_),
    .Q(\Qset[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12617_ (.CLK(clknet_leaf_35_clk),
    .D(_00067_),
    .Q(\Qset[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12618_ (.CLK(clknet_leaf_34_clk),
    .D(_00068_),
    .Q(\Qset[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12619_ (.CLK(clknet_leaf_28_clk),
    .D(_00069_),
    .Q(\Qset[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12620_ (.CLK(clknet_leaf_27_clk),
    .D(_00070_),
    .Q(\Qset[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12621_ (.CLK(clknet_leaf_27_clk),
    .D(_00071_),
    .Q(\Qset[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12622_ (.CLK(clknet_leaf_1_clk),
    .D(_00072_),
    .Q(_00002_));
 sky130_fd_sc_hd__dfxtp_2 _12623_ (.CLK(clknet_leaf_51_clk),
    .D(_00073_),
    .Q(_00003_));
 sky130_fd_sc_hd__dfxtp_1 _12624_ (.CLK(clknet_leaf_53_clk),
    .D(_00074_),
    .Q(\Oset[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12625_ (.CLK(clknet_leaf_45_clk),
    .D(_00075_),
    .Q(\Oset[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12626_ (.CLK(clknet_leaf_45_clk),
    .D(_00076_),
    .Q(\Oset[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12627_ (.CLK(clknet_3_0__leaf_clk),
    .D(_00077_),
    .Q(\Oset[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12628_ (.CLK(clknet_leaf_43_clk),
    .D(_00078_),
    .Q(\Oset[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12629_ (.CLK(clknet_leaf_45_clk),
    .D(_00079_),
    .Q(\Oset[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12630_ (.CLK(clknet_leaf_44_clk),
    .D(_00080_),
    .Q(\Oset[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12631_ (.CLK(clknet_leaf_41_clk),
    .D(_00081_),
    .Q(\Oset[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12632_ (.CLK(clknet_leaf_42_clk),
    .D(_00082_),
    .Q(\Oset[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12633_ (.CLK(clknet_leaf_40_clk),
    .D(_00083_),
    .Q(\Oset[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12634_ (.CLK(clknet_leaf_37_clk),
    .D(_00084_),
    .Q(\Oset[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12635_ (.CLK(clknet_leaf_38_clk),
    .D(_00085_),
    .Q(\Oset[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12636_ (.CLK(clknet_leaf_34_clk),
    .D(_00086_),
    .Q(\Oset[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12637_ (.CLK(clknet_leaf_28_clk),
    .D(_00087_),
    .Q(\Oset[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12638_ (.CLK(clknet_leaf_30_clk),
    .D(_00088_),
    .Q(\Oset[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12639_ (.CLK(clknet_leaf_30_clk),
    .D(_00089_),
    .Q(\Oset[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12640_ (.CLK(clknet_leaf_54_clk),
    .D(_00090_),
    .Q(_00004_));
 sky130_fd_sc_hd__dfxtp_4 _12641_ (.CLK(clknet_leaf_52_clk),
    .D(_00091_),
    .Q(_00005_));
 sky130_fd_sc_hd__dfxtp_1 _12642_ (.CLK(clknet_leaf_51_clk),
    .D(_00092_),
    .Q(_00000_));
 sky130_fd_sc_hd__dfxtp_4 _12643_ (.CLK(clknet_leaf_51_clk),
    .D(_00093_),
    .Q(_00001_));
 sky130_fd_sc_hd__dfxtp_1 _12644_ (.CLK(clknet_leaf_49_clk),
    .D(_00094_),
    .Q(\H[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12645_ (.CLK(clknet_leaf_53_clk),
    .D(_00095_),
    .Q(\H[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12646_ (.CLK(clknet_leaf_49_clk),
    .D(_00096_),
    .Q(\H[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12647_ (.CLK(clknet_leaf_46_clk),
    .D(_00097_),
    .Q(\H[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12648_ (.CLK(clknet_leaf_32_clk),
    .D(_00098_),
    .Q(\H[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12649_ (.CLK(clknet_leaf_41_clk),
    .D(_00099_),
    .Q(\H[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12650_ (.CLK(clknet_leaf_41_clk),
    .D(_00100_),
    .Q(\H[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12651_ (.CLK(clknet_leaf_32_clk),
    .D(_00101_),
    .Q(\H[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12652_ (.CLK(clknet_leaf_37_clk),
    .D(_00102_),
    .Q(\H[3][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12653_ (.CLK(clknet_leaf_40_clk),
    .D(_00103_),
    .Q(\H[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12654_ (.CLK(clknet_leaf_33_clk),
    .D(_00104_),
    .Q(\H[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12655_ (.CLK(clknet_leaf_33_clk),
    .D(_00105_),
    .Q(\H[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12656_ (.CLK(clknet_leaf_26_clk),
    .D(_00106_),
    .Q(\H[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12657_ (.CLK(clknet_leaf_26_clk),
    .D(_00107_),
    .Q(\H[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12658_ (.CLK(clknet_leaf_27_clk),
    .D(_00108_),
    .Q(\H[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12659_ (.CLK(clknet_leaf_26_clk),
    .D(_00109_),
    .Q(\H[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12660_ (.CLK(clknet_leaf_53_clk),
    .D(_00110_),
    .Q(\Oset[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12661_ (.CLK(clknet_leaf_53_clk),
    .D(_00111_),
    .Q(\Oset[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12662_ (.CLK(clknet_leaf_45_clk),
    .D(_00112_),
    .Q(\Oset[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12663_ (.CLK(clknet_3_0__leaf_clk),
    .D(_00113_),
    .Q(\Oset[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12664_ (.CLK(clknet_leaf_43_clk),
    .D(_00114_),
    .Q(\Oset[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12665_ (.CLK(clknet_leaf_45_clk),
    .D(_00115_),
    .Q(\Oset[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12666_ (.CLK(clknet_leaf_44_clk),
    .D(_00116_),
    .Q(\Oset[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12667_ (.CLK(clknet_leaf_41_clk),
    .D(_00117_),
    .Q(\Oset[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12668_ (.CLK(clknet_leaf_42_clk),
    .D(_00118_),
    .Q(\Oset[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12669_ (.CLK(clknet_leaf_40_clk),
    .D(_00119_),
    .Q(\Oset[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12670_ (.CLK(clknet_leaf_37_clk),
    .D(_00120_),
    .Q(\Oset[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12671_ (.CLK(clknet_leaf_38_clk),
    .D(_00121_),
    .Q(\Oset[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12672_ (.CLK(clknet_leaf_34_clk),
    .D(_00122_),
    .Q(\Oset[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12673_ (.CLK(clknet_leaf_28_clk),
    .D(_00123_),
    .Q(\Oset[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12674_ (.CLK(clknet_leaf_26_clk),
    .D(_00124_),
    .Q(\Oset[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12675_ (.CLK(clknet_leaf_30_clk),
    .D(_00125_),
    .Q(\Oset[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12676_ (.CLK(clknet_leaf_0_clk),
    .D(_00126_),
    .Q(\LC[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12677_ (.CLK(clknet_leaf_0_clk),
    .D(_00127_),
    .Q(\LC[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12678_ (.CLK(clknet_leaf_0_clk),
    .D(_00128_),
    .Q(\LC[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12679_ (.CLK(clknet_leaf_1_clk),
    .D(_00129_),
    .Q(\LC[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12680_ (.CLK(clknet_leaf_1_clk),
    .D(_00130_),
    .Q(\LC[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12681_ (.CLK(clknet_leaf_1_clk),
    .D(_00131_),
    .Q(\LC[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12682_ (.CLK(clknet_leaf_1_clk),
    .D(_00132_),
    .Q(\LC[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12683_ (.CLK(clknet_leaf_1_clk),
    .D(_00133_),
    .Q(\LC[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12684_ (.CLK(clknet_leaf_1_clk),
    .D(_00134_),
    .Q(\LC[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12685_ (.CLK(clknet_leaf_1_clk),
    .D(_00135_),
    .Q(\LC[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12686_ (.CLK(clknet_leaf_53_clk),
    .D(_00136_),
    .Q(\Oset[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12687_ (.CLK(clknet_leaf_53_clk),
    .D(_00137_),
    .Q(\Oset[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12688_ (.CLK(clknet_leaf_45_clk),
    .D(_00138_),
    .Q(\Oset[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12689_ (.CLK(clknet_leaf_52_clk),
    .D(_00139_),
    .Q(\Oset[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12690_ (.CLK(clknet_leaf_43_clk),
    .D(_00140_),
    .Q(\Oset[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12691_ (.CLK(clknet_leaf_45_clk),
    .D(_00141_),
    .Q(\Oset[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12692_ (.CLK(clknet_leaf_44_clk),
    .D(_00142_),
    .Q(\Oset[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12693_ (.CLK(clknet_leaf_40_clk),
    .D(_00143_),
    .Q(\Oset[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12694_ (.CLK(clknet_leaf_42_clk),
    .D(_00144_),
    .Q(\Oset[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12695_ (.CLK(clknet_leaf_40_clk),
    .D(_00145_),
    .Q(\Oset[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12696_ (.CLK(clknet_leaf_36_clk),
    .D(_00146_),
    .Q(\Oset[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12697_ (.CLK(clknet_leaf_38_clk),
    .D(_00147_),
    .Q(\Oset[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12698_ (.CLK(clknet_leaf_34_clk),
    .D(_00148_),
    .Q(\Oset[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12699_ (.CLK(clknet_leaf_29_clk),
    .D(_00149_),
    .Q(\Oset[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12700_ (.CLK(clknet_leaf_26_clk),
    .D(_00150_),
    .Q(\Oset[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12701_ (.CLK(clknet_leaf_30_clk),
    .D(_00151_),
    .Q(\Oset[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12702_ (.CLK(clknet_leaf_3_clk),
    .D(net35),
    .Q(\current_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12703_ (.CLK(clknet_leaf_3_clk),
    .D(_00008_),
    .Q(\current_state[1] ));
 sky130_fd_sc_hd__dfxtp_4 _12704_ (.CLK(clknet_leaf_3_clk),
    .D(_00009_),
    .Q(\current_state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12705_ (.CLK(clknet_leaf_5_clk),
    .D(_00013_),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_1 _12706_ (.CLK(clknet_leaf_3_clk),
    .D(_00010_),
    .Q(\current_state[4] ));
 sky130_fd_sc_hd__dfxtp_2 _12707_ (.CLK(clknet_leaf_2_clk),
    .D(_00011_),
    .Q(\current_state[5] ));
 sky130_fd_sc_hd__dfxtp_2 _12708_ (.CLK(clknet_leaf_3_clk),
    .D(_00012_),
    .Q(\current_state[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12709_ (.CLK(clknet_leaf_45_clk),
    .D(_00152_),
    .Q(\Oset[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12710_ (.CLK(clknet_leaf_53_clk),
    .D(_00153_),
    .Q(\Oset[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12711_ (.CLK(clknet_leaf_45_clk),
    .D(_00154_),
    .Q(\Oset[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12712_ (.CLK(clknet_leaf_52_clk),
    .D(_00155_),
    .Q(\Oset[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12713_ (.CLK(clknet_leaf_44_clk),
    .D(_00156_),
    .Q(\Oset[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12714_ (.CLK(clknet_leaf_45_clk),
    .D(_00157_),
    .Q(\Oset[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12715_ (.CLK(clknet_leaf_44_clk),
    .D(_00158_),
    .Q(\Oset[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12716_ (.CLK(clknet_leaf_41_clk),
    .D(_00159_),
    .Q(\Oset[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12717_ (.CLK(clknet_leaf_41_clk),
    .D(_00160_),
    .Q(\Oset[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12718_ (.CLK(clknet_leaf_40_clk),
    .D(_00161_),
    .Q(\Oset[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12719_ (.CLK(clknet_leaf_36_clk),
    .D(_00162_),
    .Q(\Oset[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12720_ (.CLK(clknet_leaf_38_clk),
    .D(_00163_),
    .Q(\Oset[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12721_ (.CLK(clknet_leaf_33_clk),
    .D(_00164_),
    .Q(\Oset[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12722_ (.CLK(clknet_leaf_28_clk),
    .D(_00165_),
    .Q(\Oset[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12723_ (.CLK(clknet_leaf_30_clk),
    .D(_00166_),
    .Q(\Oset[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12724_ (.CLK(clknet_leaf_30_clk),
    .D(_00167_),
    .Q(\Oset[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12725_ (.CLK(clknet_leaf_49_clk),
    .D(_00168_),
    .Q(\H[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12726_ (.CLK(clknet_leaf_53_clk),
    .D(_00169_),
    .Q(\H[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12727_ (.CLK(clknet_leaf_49_clk),
    .D(_00170_),
    .Q(\H[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12728_ (.CLK(clknet_leaf_44_clk),
    .D(_00171_),
    .Q(\H[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12729_ (.CLK(clknet_leaf_32_clk),
    .D(_00172_),
    .Q(\H[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12730_ (.CLK(clknet_leaf_44_clk),
    .D(_00173_),
    .Q(\H[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12731_ (.CLK(clknet_leaf_41_clk),
    .D(_00174_),
    .Q(\H[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12732_ (.CLK(clknet_leaf_37_clk),
    .D(_00175_),
    .Q(\H[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12733_ (.CLK(clknet_leaf_40_clk),
    .D(_00176_),
    .Q(\H[2][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12734_ (.CLK(clknet_leaf_40_clk),
    .D(_00177_),
    .Q(\H[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12735_ (.CLK(clknet_leaf_33_clk),
    .D(_00178_),
    .Q(\H[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12736_ (.CLK(clknet_leaf_33_clk),
    .D(_00179_),
    .Q(\H[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12737_ (.CLK(clknet_leaf_26_clk),
    .D(_00180_),
    .Q(\H[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12738_ (.CLK(clknet_leaf_25_clk),
    .D(_00181_),
    .Q(\H[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12739_ (.CLK(clknet_leaf_25_clk),
    .D(_00182_),
    .Q(\H[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12740_ (.CLK(clknet_leaf_26_clk),
    .D(_00183_),
    .Q(\H[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12741_ (.CLK(clknet_leaf_49_clk),
    .D(_00184_),
    .Q(\H[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12742_ (.CLK(clknet_leaf_53_clk),
    .D(_00185_),
    .Q(\H[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12743_ (.CLK(clknet_leaf_49_clk),
    .D(_00186_),
    .Q(\H[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12744_ (.CLK(clknet_leaf_45_clk),
    .D(_00187_),
    .Q(\H[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12745_ (.CLK(clknet_leaf_32_clk),
    .D(_00188_),
    .Q(\H[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12746_ (.CLK(clknet_leaf_41_clk),
    .D(_00189_),
    .Q(\H[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12747_ (.CLK(clknet_leaf_41_clk),
    .D(_00190_),
    .Q(\H[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12748_ (.CLK(clknet_leaf_37_clk),
    .D(_00191_),
    .Q(\H[1][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12749_ (.CLK(clknet_leaf_40_clk),
    .D(_00192_),
    .Q(\H[1][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12750_ (.CLK(clknet_leaf_40_clk),
    .D(_00193_),
    .Q(\H[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12751_ (.CLK(clknet_leaf_33_clk),
    .D(_00194_),
    .Q(\H[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12752_ (.CLK(clknet_leaf_33_clk),
    .D(_00195_),
    .Q(\H[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12753_ (.CLK(clknet_leaf_26_clk),
    .D(_00196_),
    .Q(\H[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12754_ (.CLK(clknet_leaf_26_clk),
    .D(_00197_),
    .Q(\H[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12755_ (.CLK(clknet_leaf_26_clk),
    .D(_00198_),
    .Q(\H[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12756_ (.CLK(clknet_leaf_30_clk),
    .D(_00199_),
    .Q(\H[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12757_ (.CLK(clknet_leaf_49_clk),
    .D(_00200_),
    .Q(\H[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12758_ (.CLK(clknet_leaf_53_clk),
    .D(_00201_),
    .Q(\H[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12759_ (.CLK(clknet_leaf_49_clk),
    .D(_00202_),
    .Q(\H[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12760_ (.CLK(clknet_leaf_45_clk),
    .D(_00203_),
    .Q(\H[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12761_ (.CLK(clknet_leaf_32_clk),
    .D(_00204_),
    .Q(\H[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12762_ (.CLK(clknet_leaf_43_clk),
    .D(_00205_),
    .Q(\H[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12763_ (.CLK(clknet_leaf_41_clk),
    .D(_00206_),
    .Q(\H[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12764_ (.CLK(clknet_leaf_37_clk),
    .D(_00207_),
    .Q(\H[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12765_ (.CLK(clknet_leaf_40_clk),
    .D(_00208_),
    .Q(\H[0][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12766_ (.CLK(clknet_leaf_40_clk),
    .D(_00209_),
    .Q(\H[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12767_ (.CLK(clknet_leaf_33_clk),
    .D(_00210_),
    .Q(\H[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12768_ (.CLK(clknet_leaf_33_clk),
    .D(_00211_),
    .Q(\H[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12769_ (.CLK(clknet_leaf_26_clk),
    .D(_00212_),
    .Q(\H[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12770_ (.CLK(clknet_leaf_26_clk),
    .D(_00213_),
    .Q(\H[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12771_ (.CLK(clknet_leaf_26_clk),
    .D(_00214_),
    .Q(\H[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12772_ (.CLK(clknet_leaf_26_clk),
    .D(_00215_),
    .Q(\H[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12773_ (.CLK(clknet_leaf_27_clk),
    .D(_00216_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_1 _12774_ (.CLK(clknet_leaf_28_clk),
    .D(_00217_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _12775_ (.CLK(clknet_leaf_27_clk),
    .D(_00218_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _12776_ (.CLK(clknet_leaf_27_clk),
    .D(_00219_),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _12777_ (.CLK(clknet_leaf_25_clk),
    .D(_00220_),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_1 _12778_ (.CLK(clknet_leaf_25_clk),
    .D(_00221_),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_1 _12779_ (.CLK(clknet_leaf_24_clk),
    .D(_00222_),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_1 _12780_ (.CLK(clknet_leaf_24_clk),
    .D(_00223_),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_1 _12781_ (.CLK(clknet_leaf_24_clk),
    .D(_00224_),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_1 _12782_ (.CLK(clknet_leaf_27_clk),
    .D(_00225_),
    .Q(net47));
 sky130_fd_sc_hd__dfxtp_4 _12783_ (.CLK(clknet_leaf_28_clk),
    .D(_00226_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _12784_ (.CLK(clknet_leaf_2_clk),
    .D(_00227_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _12785_ (.CLK(clknet_leaf_54_clk),
    .D(_00228_),
    .Q(net48));
 sky130_fd_sc_hd__dfxtp_1 _12786_ (.CLK(clknet_leaf_54_clk),
    .D(_00229_),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_1 _12787_ (.CLK(clknet_leaf_54_clk),
    .D(_00230_),
    .Q(net56));
 sky130_fd_sc_hd__dfxtp_1 _12788_ (.CLK(clknet_leaf_54_clk),
    .D(_00231_),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_1 _12789_ (.CLK(clknet_leaf_53_clk),
    .D(_00232_),
    .Q(net58));
 sky130_fd_sc_hd__dfxtp_1 _12790_ (.CLK(clknet_leaf_45_clk),
    .D(_00233_),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_1 _12791_ (.CLK(clknet_leaf_45_clk),
    .D(_00234_),
    .Q(net60));
 sky130_fd_sc_hd__dfxtp_1 _12792_ (.CLK(clknet_leaf_45_clk),
    .D(_00235_),
    .Q(net61));
 sky130_fd_sc_hd__dfxtp_1 _12793_ (.CLK(clknet_leaf_44_clk),
    .D(_00236_),
    .Q(net62));
 sky130_fd_sc_hd__dfxtp_1 _12794_ (.CLK(clknet_leaf_44_clk),
    .D(_00237_),
    .Q(net63));
 sky130_fd_sc_hd__dfxtp_1 _12795_ (.CLK(clknet_leaf_44_clk),
    .D(_00238_),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_1 _12796_ (.CLK(clknet_leaf_41_clk),
    .D(_00239_),
    .Q(net50));
 sky130_fd_sc_hd__dfxtp_1 _12797_ (.CLK(clknet_leaf_40_clk),
    .D(_00240_),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_1 _12798_ (.CLK(clknet_leaf_40_clk),
    .D(_00241_),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_1 _12799_ (.CLK(clknet_leaf_40_clk),
    .D(_00242_),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_1 _12800_ (.CLK(clknet_leaf_39_clk),
    .D(_00243_),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_1 _12801_ (.CLK(clknet_leaf_10_clk),
    .D(_00244_),
    .Q(\result_reg_add[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12802_ (.CLK(clknet_leaf_9_clk),
    .D(_00245_),
    .Q(\result_reg_add[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12803_ (.CLK(clknet_leaf_11_clk),
    .D(_00246_),
    .Q(\result_reg_add[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12804_ (.CLK(clknet_leaf_11_clk),
    .D(_00247_),
    .Q(\result_reg_add[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12805_ (.CLK(clknet_leaf_11_clk),
    .D(_00248_),
    .Q(\result_reg_add[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12806_ (.CLK(clknet_leaf_11_clk),
    .D(_00249_),
    .Q(\result_reg_add[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12807_ (.CLK(clknet_leaf_11_clk),
    .D(_00250_),
    .Q(\result_reg_add[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12808_ (.CLK(clknet_leaf_12_clk),
    .D(_00251_),
    .Q(\result_reg_add[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12809_ (.CLK(clknet_leaf_10_clk),
    .D(_00252_),
    .Q(\result_reg_add[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12810_ (.CLK(clknet_leaf_12_clk),
    .D(_00253_),
    .Q(\result_reg_add[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12811_ (.CLK(clknet_leaf_12_clk),
    .D(_00254_),
    .Q(\result_reg_add[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12812_ (.CLK(clknet_leaf_10_clk),
    .D(_00255_),
    .Q(\result_reg_add[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12813_ (.CLK(clknet_leaf_9_clk),
    .D(_00256_),
    .Q(\result_reg_add[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12814_ (.CLK(clknet_leaf_9_clk),
    .D(_00257_),
    .Q(\result_reg_add[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12815_ (.CLK(clknet_leaf_10_clk),
    .D(_00258_),
    .Q(\result_reg_add[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12816_ (.CLK(clknet_leaf_10_clk),
    .D(_00259_),
    .Q(\result_reg_add[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12817_ (.CLK(clknet_leaf_10_clk),
    .D(_00260_),
    .Q(\result_reg_sub[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12818_ (.CLK(clknet_leaf_10_clk),
    .D(_00261_),
    .Q(\result_reg_sub[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12819_ (.CLK(clknet_leaf_11_clk),
    .D(_00262_),
    .Q(\result_reg_sub[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12820_ (.CLK(clknet_leaf_11_clk),
    .D(_00263_),
    .Q(\result_reg_sub[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12821_ (.CLK(clknet_leaf_11_clk),
    .D(_00264_),
    .Q(\result_reg_sub[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12822_ (.CLK(clknet_leaf_10_clk),
    .D(_00265_),
    .Q(\result_reg_sub[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12823_ (.CLK(clknet_leaf_11_clk),
    .D(_00266_),
    .Q(\result_reg_sub[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12824_ (.CLK(clknet_leaf_12_clk),
    .D(_00267_),
    .Q(\result_reg_sub[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12825_ (.CLK(clknet_leaf_10_clk),
    .D(_00268_),
    .Q(\result_reg_sub[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12826_ (.CLK(clknet_leaf_12_clk),
    .D(_00269_),
    .Q(\result_reg_sub[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12827_ (.CLK(clknet_leaf_12_clk),
    .D(_00270_),
    .Q(\result_reg_sub[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12828_ (.CLK(clknet_leaf_10_clk),
    .D(_00271_),
    .Q(\result_reg_sub[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12829_ (.CLK(clknet_leaf_9_clk),
    .D(_00272_),
    .Q(\result_reg_sub[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12830_ (.CLK(clknet_leaf_8_clk),
    .D(_00273_),
    .Q(\result_reg_sub[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12831_ (.CLK(clknet_leaf_9_clk),
    .D(_00274_),
    .Q(\result_reg_sub[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12832_ (.CLK(clknet_leaf_10_clk),
    .D(_00275_),
    .Q(\result_reg_sub[15] ));
 sky130_fd_sc_hd__dfxtp_2 _12833_ (.CLK(clknet_leaf_2_clk),
    .D(_00276_),
    .Q(\result_reg_mul[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12834_ (.CLK(clknet_leaf_7_clk),
    .D(_00277_),
    .Q(\result_reg_mul[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12835_ (.CLK(clknet_leaf_8_clk),
    .D(_00278_),
    .Q(\result_reg_mul[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12836_ (.CLK(clknet_leaf_7_clk),
    .D(_00279_),
    .Q(\result_reg_mul[3] ));
 sky130_fd_sc_hd__dfxtp_2 _12837_ (.CLK(clknet_leaf_56_clk),
    .D(_00280_),
    .Q(\result_reg_mul[4] ));
 sky130_fd_sc_hd__dfxtp_2 _12838_ (.CLK(clknet_leaf_4_clk),
    .D(_00281_),
    .Q(\result_reg_mul[5] ));
 sky130_fd_sc_hd__dfxtp_2 _12839_ (.CLK(clknet_leaf_0_clk),
    .D(_00282_),
    .Q(\result_reg_mul[6] ));
 sky130_fd_sc_hd__dfxtp_2 _12840_ (.CLK(clknet_leaf_56_clk),
    .D(_00283_),
    .Q(\result_reg_mul[7] ));
 sky130_fd_sc_hd__dfxtp_2 _12841_ (.CLK(clknet_leaf_56_clk),
    .D(_00284_),
    .Q(\result_reg_mul[8] ));
 sky130_fd_sc_hd__dfxtp_2 _12842_ (.CLK(clknet_leaf_56_clk),
    .D(_00285_),
    .Q(\result_reg_mul[9] ));
 sky130_fd_sc_hd__dfxtp_2 _12843_ (.CLK(clknet_leaf_56_clk),
    .D(_00286_),
    .Q(\result_reg_mul[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12844_ (.CLK(clknet_leaf_8_clk),
    .D(_00287_),
    .Q(\result_reg_mul[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12845_ (.CLK(clknet_leaf_4_clk),
    .D(_00288_),
    .Q(\result_reg_mul[12] ));
 sky130_fd_sc_hd__dfxtp_2 _12846_ (.CLK(clknet_leaf_4_clk),
    .D(_00289_),
    .Q(\result_reg_mul[13] ));
 sky130_fd_sc_hd__dfxtp_2 _12847_ (.CLK(clknet_leaf_5_clk),
    .D(_00290_),
    .Q(\result_reg_mul[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12848_ (.CLK(clknet_leaf_7_clk),
    .D(_00291_),
    .Q(\result_reg_mul[15] ));
 sky130_fd_sc_hd__dfxtp_2 _12849_ (.CLK(clknet_leaf_10_clk),
    .D(_00292_),
    .Q(\result_reg_mac[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12850_ (.CLK(clknet_leaf_20_clk),
    .D(_00293_),
    .Q(\result_reg_mac[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12851_ (.CLK(clknet_leaf_18_clk),
    .D(_00294_),
    .Q(\result_reg_mac[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12852_ (.CLK(clknet_leaf_18_clk),
    .D(_00295_),
    .Q(\result_reg_mac[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12853_ (.CLK(clknet_leaf_18_clk),
    .D(_00296_),
    .Q(\result_reg_mac[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12854_ (.CLK(clknet_leaf_18_clk),
    .D(_00297_),
    .Q(\result_reg_mac[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12855_ (.CLK(clknet_leaf_18_clk),
    .D(_00298_),
    .Q(\result_reg_mac[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12856_ (.CLK(clknet_leaf_18_clk),
    .D(_00299_),
    .Q(\result_reg_mac[7] ));
 sky130_fd_sc_hd__dfxtp_2 _12857_ (.CLK(clknet_leaf_10_clk),
    .D(_00300_),
    .Q(\result_reg_mac[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12858_ (.CLK(clknet_leaf_18_clk),
    .D(_00301_),
    .Q(\result_reg_mac[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12859_ (.CLK(clknet_leaf_18_clk),
    .D(_00302_),
    .Q(\result_reg_mac[10] ));
 sky130_fd_sc_hd__dfxtp_2 _12860_ (.CLK(clknet_leaf_10_clk),
    .D(_00303_),
    .Q(\result_reg_mac[11] ));
 sky130_fd_sc_hd__dfxtp_2 _12861_ (.CLK(clknet_leaf_8_clk),
    .D(_00304_),
    .Q(\result_reg_mac[12] ));
 sky130_fd_sc_hd__dfxtp_2 _12862_ (.CLK(clknet_leaf_9_clk),
    .D(_00305_),
    .Q(\result_reg_mac[13] ));
 sky130_fd_sc_hd__dfxtp_2 _12863_ (.CLK(clknet_leaf_10_clk),
    .D(_00306_),
    .Q(\result_reg_mac[14] ));
 sky130_fd_sc_hd__dfxtp_2 _12864_ (.CLK(clknet_leaf_10_clk),
    .D(_00307_),
    .Q(\result_reg_mac[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12865_ (.CLK(clknet_leaf_20_clk),
    .D(_00308_),
    .Q(\result_reg_Lshift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12866_ (.CLK(clknet_leaf_24_clk),
    .D(_00309_),
    .Q(\result_reg_Lshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12867_ (.CLK(clknet_leaf_23_clk),
    .D(_00310_),
    .Q(\result_reg_Lshift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12868_ (.CLK(clknet_leaf_23_clk),
    .D(_00311_),
    .Q(\result_reg_Lshift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12869_ (.CLK(clknet_leaf_19_clk),
    .D(_00312_),
    .Q(\result_reg_Lshift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12870_ (.CLK(clknet_leaf_23_clk),
    .D(_00313_),
    .Q(\result_reg_Lshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12871_ (.CLK(clknet_leaf_23_clk),
    .D(_00314_),
    .Q(\result_reg_Lshift[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12872_ (.CLK(clknet_leaf_22_clk),
    .D(_00315_),
    .Q(\result_reg_Lshift[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12873_ (.CLK(clknet_leaf_24_clk),
    .D(_00316_),
    .Q(\result_reg_Lshift[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12874_ (.CLK(clknet_leaf_24_clk),
    .D(_00317_),
    .Q(\result_reg_Lshift[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12875_ (.CLK(clknet_leaf_24_clk),
    .D(_00318_),
    .Q(\result_reg_Lshift[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12876_ (.CLK(clknet_leaf_24_clk),
    .D(_00319_),
    .Q(\result_reg_Lshift[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12877_ (.CLK(clknet_leaf_25_clk),
    .D(_00320_),
    .Q(\result_reg_Lshift[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12878_ (.CLK(clknet_leaf_25_clk),
    .D(_00321_),
    .Q(\result_reg_Lshift[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12879_ (.CLK(clknet_leaf_24_clk),
    .D(_00322_),
    .Q(\result_reg_Lshift[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12880_ (.CLK(clknet_leaf_20_clk),
    .D(_00323_),
    .Q(\result_reg_Lshift[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12881_ (.CLK(clknet_leaf_21_clk),
    .D(_00324_),
    .Q(\result_reg_Rshift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12882_ (.CLK(clknet_leaf_24_clk),
    .D(_00325_),
    .Q(\result_reg_Rshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12883_ (.CLK(clknet_leaf_23_clk),
    .D(_00326_),
    .Q(\result_reg_Rshift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12884_ (.CLK(clknet_leaf_23_clk),
    .D(_00327_),
    .Q(\result_reg_Rshift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12885_ (.CLK(clknet_leaf_19_clk),
    .D(_00328_),
    .Q(\result_reg_Rshift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12886_ (.CLK(clknet_leaf_23_clk),
    .D(_00329_),
    .Q(\result_reg_Rshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12887_ (.CLK(clknet_leaf_23_clk),
    .D(_00330_),
    .Q(\result_reg_Rshift[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12888_ (.CLK(clknet_leaf_22_clk),
    .D(_00331_),
    .Q(\result_reg_Rshift[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12889_ (.CLK(clknet_leaf_24_clk),
    .D(_00332_),
    .Q(\result_reg_Rshift[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12890_ (.CLK(clknet_leaf_23_clk),
    .D(_00333_),
    .Q(\result_reg_Rshift[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12891_ (.CLK(clknet_leaf_24_clk),
    .D(_00334_),
    .Q(\result_reg_Rshift[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12892_ (.CLK(clknet_leaf_24_clk),
    .D(_00335_),
    .Q(\result_reg_Rshift[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12893_ (.CLK(clknet_leaf_24_clk),
    .D(_00336_),
    .Q(\result_reg_Rshift[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12894_ (.CLK(clknet_leaf_24_clk),
    .D(_00337_),
    .Q(\result_reg_Rshift[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12895_ (.CLK(clknet_leaf_24_clk),
    .D(_00338_),
    .Q(\result_reg_Rshift[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12896_ (.CLK(clknet_leaf_21_clk),
    .D(_00339_),
    .Q(\result_reg_Rshift[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12897_ (.CLK(clknet_leaf_16_clk),
    .D(_00340_),
    .Q(\result_reg_and[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12898_ (.CLK(clknet_leaf_14_clk),
    .D(_00341_),
    .Q(\result_reg_and[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12899_ (.CLK(clknet_leaf_15_clk),
    .D(_00342_),
    .Q(\result_reg_and[2] ));
 sky130_fd_sc_hd__dfxtp_2 _12900_ (.CLK(clknet_leaf_15_clk),
    .D(_00343_),
    .Q(\result_reg_and[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12901_ (.CLK(clknet_leaf_16_clk),
    .D(_00344_),
    .Q(\result_reg_and[4] ));
 sky130_fd_sc_hd__dfxtp_2 _12902_ (.CLK(clknet_leaf_15_clk),
    .D(_00345_),
    .Q(\result_reg_and[5] ));
 sky130_fd_sc_hd__dfxtp_2 _12903_ (.CLK(clknet_leaf_16_clk),
    .D(_00346_),
    .Q(\result_reg_and[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12904_ (.CLK(clknet_leaf_16_clk),
    .D(_00347_),
    .Q(\result_reg_and[7] ));
 sky130_fd_sc_hd__dfxtp_2 _12905_ (.CLK(clknet_leaf_31_clk),
    .D(_00348_),
    .Q(\result_reg_and[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12906_ (.CLK(clknet_leaf_17_clk),
    .D(_00349_),
    .Q(\result_reg_and[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12907_ (.CLK(clknet_leaf_16_clk),
    .D(_00350_),
    .Q(\result_reg_and[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12908_ (.CLK(clknet_leaf_16_clk),
    .D(_00351_),
    .Q(\result_reg_and[11] ));
 sky130_fd_sc_hd__dfxtp_2 _12909_ (.CLK(clknet_leaf_31_clk),
    .D(_00352_),
    .Q(\result_reg_and[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12910_ (.CLK(clknet_leaf_16_clk),
    .D(_00353_),
    .Q(\result_reg_and[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12911_ (.CLK(clknet_leaf_17_clk),
    .D(_00354_),
    .Q(\result_reg_and[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12912_ (.CLK(clknet_leaf_16_clk),
    .D(_00355_),
    .Q(\result_reg_and[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12913_ (.CLK(clknet_leaf_15_clk),
    .D(_00356_),
    .Q(\result_reg_or[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12914_ (.CLK(clknet_leaf_15_clk),
    .D(_00357_),
    .Q(\result_reg_or[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12915_ (.CLK(clknet_leaf_15_clk),
    .D(_00358_),
    .Q(\result_reg_or[2] ));
 sky130_fd_sc_hd__dfxtp_2 _12916_ (.CLK(clknet_leaf_15_clk),
    .D(_00359_),
    .Q(\result_reg_or[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12917_ (.CLK(clknet_leaf_17_clk),
    .D(_00360_),
    .Q(\result_reg_or[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12918_ (.CLK(clknet_leaf_16_clk),
    .D(_00361_),
    .Q(\result_reg_or[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12919_ (.CLK(clknet_leaf_31_clk),
    .D(_00362_),
    .Q(\result_reg_or[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12920_ (.CLK(clknet_leaf_16_clk),
    .D(_00363_),
    .Q(\result_reg_or[7] ));
 sky130_fd_sc_hd__dfxtp_2 _12921_ (.CLK(clknet_leaf_31_clk),
    .D(_00364_),
    .Q(\result_reg_or[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12922_ (.CLK(clknet_leaf_17_clk),
    .D(_00365_),
    .Q(\result_reg_or[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12923_ (.CLK(clknet_leaf_17_clk),
    .D(_00366_),
    .Q(\result_reg_or[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12924_ (.CLK(clknet_leaf_17_clk),
    .D(_00367_),
    .Q(\result_reg_or[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12925_ (.CLK(clknet_leaf_21_clk),
    .D(_00368_),
    .Q(\result_reg_or[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12926_ (.CLK(clknet_leaf_16_clk),
    .D(_00369_),
    .Q(\result_reg_or[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12927_ (.CLK(clknet_leaf_30_clk),
    .D(_00370_),
    .Q(\result_reg_or[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12928_ (.CLK(clknet_leaf_16_clk),
    .D(_00371_),
    .Q(\result_reg_or[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12929_ (.CLK(clknet_leaf_19_clk),
    .D(_00372_),
    .Q(\result_reg_not[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12930_ (.CLK(clknet_leaf_19_clk),
    .D(_00373_),
    .Q(\result_reg_not[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12931_ (.CLK(clknet_leaf_22_clk),
    .D(_00374_),
    .Q(\result_reg_not[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12932_ (.CLK(clknet_leaf_22_clk),
    .D(_00375_),
    .Q(\result_reg_not[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12933_ (.CLK(clknet_leaf_19_clk),
    .D(_00376_),
    .Q(\result_reg_not[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12934_ (.CLK(clknet_leaf_22_clk),
    .D(_00377_),
    .Q(\result_reg_not[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12935_ (.CLK(clknet_leaf_22_clk),
    .D(_00378_),
    .Q(\result_reg_not[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12936_ (.CLK(clknet_leaf_22_clk),
    .D(_00379_),
    .Q(\result_reg_not[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12937_ (.CLK(clknet_leaf_22_clk),
    .D(_00380_),
    .Q(\result_reg_not[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12938_ (.CLK(clknet_leaf_22_clk),
    .D(_00381_),
    .Q(\result_reg_not[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12939_ (.CLK(clknet_leaf_22_clk),
    .D(_00382_),
    .Q(\result_reg_not[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12940_ (.CLK(clknet_leaf_21_clk),
    .D(_00383_),
    .Q(\result_reg_not[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12941_ (.CLK(clknet_leaf_26_clk),
    .D(_00384_),
    .Q(\result_reg_not[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12942_ (.CLK(clknet_leaf_26_clk),
    .D(_00385_),
    .Q(\result_reg_not[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12943_ (.CLK(clknet_leaf_26_clk),
    .D(_00386_),
    .Q(\result_reg_not[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12944_ (.CLK(clknet_leaf_21_clk),
    .D(_00387_),
    .Q(\result_reg_not[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12945_ (.CLK(clknet_leaf_14_clk),
    .D(_00388_),
    .Q(\result_reg_set[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12946_ (.CLK(clknet_leaf_15_clk),
    .D(_00389_),
    .Q(\result_reg_set[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12947_ (.CLK(clknet_leaf_15_clk),
    .D(_00390_),
    .Q(\result_reg_set[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12948_ (.CLK(clknet_leaf_14_clk),
    .D(_00391_),
    .Q(\result_reg_set[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12949_ (.CLK(clknet_leaf_15_clk),
    .D(_00392_),
    .Q(\result_reg_set[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12950_ (.CLK(clknet_leaf_1_clk),
    .D(_00393_),
    .Q(\result_reg_set[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12951_ (.CLK(clknet_leaf_15_clk),
    .D(_00394_),
    .Q(\result_reg_set[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12952_ (.CLK(clknet_leaf_15_clk),
    .D(_00395_),
    .Q(\result_reg_set[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12953_ (.CLK(clknet_3_5__leaf_clk),
    .D(_00396_),
    .Q(\result_reg_set[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12954_ (.CLK(clknet_leaf_15_clk),
    .D(_00397_),
    .Q(\result_reg_set[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12955_ (.CLK(clknet_leaf_15_clk),
    .D(_00398_),
    .Q(\result_reg_set[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12956_ (.CLK(clknet_leaf_14_clk),
    .D(_00399_),
    .Q(\result_reg_set[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12957_ (.CLK(clknet_leaf_1_clk),
    .D(_00400_),
    .Q(\result_reg_set[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12958_ (.CLK(clknet_leaf_1_clk),
    .D(_00401_),
    .Q(\result_reg_set[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12959_ (.CLK(clknet_leaf_2_clk),
    .D(_00402_),
    .Q(\result_reg_set[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12960_ (.CLK(clknet_leaf_2_clk),
    .D(_00403_),
    .Q(\result_reg_set[15] ));
 sky130_fd_sc_hd__dfxtp_4 _12961_ (.CLK(clknet_leaf_54_clk),
    .D(_00404_),
    .Q(\R3[1] ));
 sky130_fd_sc_hd__dfxtp_4 _12962_ (.CLK(clknet_leaf_52_clk),
    .D(_00405_),
    .Q(\R2[1] ));
 sky130_fd_sc_hd__dfxtp_4 _12963_ (.CLK(clknet_3_1__leaf_clk),
    .D(_00406_),
    .Q(\R1[1] ));
 sky130_fd_sc_hd__dfxtp_4 _12964_ (.CLK(clknet_leaf_6_clk),
    .D(_00407_),
    .Q(\im_reg[6] ));
 sky130_fd_sc_hd__dfxtp_4 _12965_ (.CLK(clknet_leaf_6_clk),
    .D(_00408_),
    .Q(\im_reg[7] ));
 sky130_fd_sc_hd__dfxtp_4 _12966_ (.CLK(clknet_leaf_6_clk),
    .D(_00409_),
    .Q(\im_reg[8] ));
 sky130_fd_sc_hd__dfxtp_4 _12967_ (.CLK(clknet_leaf_6_clk),
    .D(_00410_),
    .Q(\im_reg[9] ));
 sky130_fd_sc_hd__dfxtp_2 _12968_ (.CLK(clknet_leaf_7_clk),
    .D(_00411_),
    .Q(CMD_addition));
 sky130_fd_sc_hd__dfxtp_1 _12969_ (.CLK(clknet_leaf_7_clk),
    .D(_00412_),
    .Q(CMD_multiplication));
 sky130_fd_sc_hd__dfxtp_1 _12970_ (.CLK(clknet_leaf_3_clk),
    .D(_00413_),
    .Q(\Add.sub ));
 sky130_fd_sc_hd__dfxtp_1 _12971_ (.CLK(clknet_leaf_1_clk),
    .D(_00414_),
    .Q(CMD_mul_accumulation));
 sky130_fd_sc_hd__dfxtp_2 _12972_ (.CLK(clknet_leaf_7_clk),
    .D(_00415_),
    .Q(CMD_logic_shift_right));
 sky130_fd_sc_hd__dfxtp_2 _12973_ (.CLK(clknet_leaf_3_clk),
    .D(_00416_),
    .Q(\shift.left ));
 sky130_fd_sc_hd__dfxtp_1 _12974_ (.CLK(clknet_leaf_3_clk),
    .D(_00417_),
    .Q(CMD_and));
 sky130_fd_sc_hd__dfxtp_1 _12975_ (.CLK(clknet_leaf_7_clk),
    .D(_00418_),
    .Q(CMD_or));
 sky130_fd_sc_hd__dfxtp_2 _12976_ (.CLK(clknet_leaf_7_clk),
    .D(_00419_),
    .Q(CMD_not));
 sky130_fd_sc_hd__dfxtp_1 _12977_ (.CLK(clknet_leaf_7_clk),
    .D(_00420_),
    .Q(CMD_load));
 sky130_fd_sc_hd__dfxtp_1 _12978_ (.CLK(clknet_leaf_7_clk),
    .D(_00421_),
    .Q(CMD_store));
 sky130_fd_sc_hd__dfxtp_1 _12979_ (.CLK(clknet_leaf_2_clk),
    .D(_00422_),
    .Q(CMD_set));
 sky130_fd_sc_hd__dfxtp_1 _12980_ (.CLK(clknet_leaf_3_clk),
    .D(_00423_),
    .Q(CMD_loopjump));
 sky130_fd_sc_hd__dfxtp_1 _12981_ (.CLK(clknet_leaf_2_clk),
    .D(_00424_),
    .Q(CMD_setloop));
 sky130_fd_sc_hd__dfxtp_2 _12982_ (.CLK(clknet_leaf_3_clk),
    .D(_00425_),
    .Q(\shift.H ));
 sky130_fd_sc_hd__dfxtp_4 _12983_ (.CLK(clknet_leaf_7_clk),
    .D(_00426_),
    .Q(Hreg2));
 sky130_fd_sc_hd__dfxtp_2 _12984_ (.CLK(clknet_leaf_2_clk),
    .D(_00427_),
    .Q(Hreg3));
 sky130_fd_sc_hd__dfxtp_1 _12985_ (.CLK(clknet_leaf_7_clk),
    .D(_00428_),
    .Q(Him));
 sky130_fd_sc_hd__dfxtp_1 _12986_ (.CLK(clknet_leaf_5_clk),
    .D(_00429_),
    .Q(\shift.O ));
 sky130_fd_sc_hd__dfxtp_4 _12987_ (.CLK(clknet_leaf_6_clk),
    .D(_00430_),
    .Q(Oreg2));
 sky130_fd_sc_hd__dfxtp_2 _12988_ (.CLK(clknet_leaf_0_clk),
    .D(_00431_),
    .Q(Oreg3));
 sky130_fd_sc_hd__dfxtp_1 _12989_ (.CLK(clknet_leaf_7_clk),
    .D(_00432_),
    .Q(Oim));
 sky130_fd_sc_hd__dfxtp_1 _12990_ (.CLK(clknet_leaf_0_clk),
    .D(_00433_),
    .Q(\shift.Q ));
 sky130_fd_sc_hd__dfxtp_1 _12991_ (.CLK(clknet_leaf_6_clk),
    .D(_00434_),
    .Q(Qreg2));
 sky130_fd_sc_hd__dfxtp_1 _12992_ (.CLK(clknet_leaf_2_clk),
    .D(_00435_),
    .Q(Qreg3));
 sky130_fd_sc_hd__dfxtp_1 _12993_ (.CLK(clknet_leaf_7_clk),
    .D(_00436_),
    .Q(Qim));
 sky130_fd_sc_hd__dfxtp_2 _12994_ (.CLK(clknet_leaf_7_clk),
    .D(_00437_),
    .Q(\R0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12995_ (.CLK(clknet_leaf_15_clk),
    .D(_00438_),
    .Q(\R0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12996_ (.CLK(clknet_leaf_0_clk),
    .D(_00439_),
    .Q(\R1[0] ));
 sky130_fd_sc_hd__dfxtp_4 _12997_ (.CLK(clknet_3_0__leaf_clk),
    .D(_00440_),
    .Q(\R2[0] ));
 sky130_fd_sc_hd__dfxtp_4 _12998_ (.CLK(clknet_leaf_54_clk),
    .D(_00441_),
    .Q(\R3[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12999_ (.CLK(clknet_leaf_39_clk),
    .D(_00442_),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_1 _13000_ (.CLK(clknet_leaf_39_clk),
    .D(_00443_),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_1 _13001_ (.CLK(clknet_leaf_39_clk),
    .D(_00444_),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_1 _13002_ (.CLK(clknet_leaf_38_clk),
    .D(_00445_),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_1 _13003_ (.CLK(clknet_leaf_38_clk),
    .D(_00446_),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_1 _13004_ (.CLK(clknet_leaf_36_clk),
    .D(_00447_),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_1 _13005_ (.CLK(clknet_leaf_35_clk),
    .D(_00448_),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_1 _13006_ (.CLK(clknet_leaf_35_clk),
    .D(_00449_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_1 _13007_ (.CLK(clknet_leaf_35_clk),
    .D(_00450_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_1 _13008_ (.CLK(clknet_leaf_34_clk),
    .D(_00451_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_1 _13009_ (.CLK(clknet_leaf_49_clk),
    .D(_00452_),
    .Q(\Qset[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13010_ (.CLK(clknet_leaf_46_clk),
    .D(_00453_),
    .Q(\Qset[3][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13011_ (.CLK(clknet_leaf_46_clk),
    .D(_00454_),
    .Q(\Qset[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13012_ (.CLK(clknet_leaf_48_clk),
    .D(_00455_),
    .Q(\Qset[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13013_ (.CLK(clknet_leaf_48_clk),
    .D(_00456_),
    .Q(\Qset[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13014_ (.CLK(clknet_leaf_46_clk),
    .D(_00457_),
    .Q(\Qset[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13015_ (.CLK(clknet_leaf_44_clk),
    .D(_00458_),
    .Q(\Qset[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13016_ (.CLK(clknet_leaf_43_clk),
    .D(_00459_),
    .Q(\Qset[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13017_ (.CLK(clknet_leaf_39_clk),
    .D(_00460_),
    .Q(\Qset[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13018_ (.CLK(clknet_leaf_39_clk),
    .D(_00461_),
    .Q(\Qset[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13019_ (.CLK(clknet_leaf_35_clk),
    .D(_00462_),
    .Q(\Qset[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13020_ (.CLK(clknet_leaf_35_clk),
    .D(_00463_),
    .Q(\Qset[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13021_ (.CLK(clknet_leaf_29_clk),
    .D(_00464_),
    .Q(\Qset[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13022_ (.CLK(clknet_leaf_28_clk),
    .D(_00465_),
    .Q(\Qset[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13023_ (.CLK(clknet_leaf_25_clk),
    .D(_00466_),
    .Q(\Qset[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13024_ (.CLK(clknet_leaf_25_clk),
    .D(_00467_),
    .Q(\Qset[3][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13025_ (.CLK(clknet_leaf_52_clk),
    .D(_00468_),
    .Q(_00006_));
 sky130_fd_sc_hd__dfxtp_2 _13026_ (.CLK(clknet_leaf_54_clk),
    .D(_00469_),
    .Q(_00007_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_38_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_39_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_40_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_41_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_42_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_43_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_44_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_45_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_46_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_48_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_49_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_51_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_52_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_53_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_54_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_56_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(data_in[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(data_in[3]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(data_in[4]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(data_in[5]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(data_in[6]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(data_in[7]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(data_in[8]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(data_in[9]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(instruction_in[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(instruction_in[10]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(instruction_in[11]),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(data_in[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input20 (.A(instruction_in[12]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(instruction_in[13]),
    .X(net21));
 sky130_fd_sc_hd__buf_2 input22 (.A(instruction_in[14]),
    .X(net22));
 sky130_fd_sc_hd__buf_2 input23 (.A(instruction_in[15]),
    .X(net23));
 sky130_fd_sc_hd__buf_2 input24 (.A(instruction_in[16]),
    .X(net24));
 sky130_fd_sc_hd__buf_2 input25 (.A(instruction_in[17]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(instruction_in[1]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(instruction_in[2]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(instruction_in[3]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(instruction_in[4]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(data_in[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input30 (.A(instruction_in[5]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(instruction_in[6]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(instruction_in[7]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(instruction_in[8]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(instruction_in[9]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(rst),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(data_in[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(data_in[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(data_in[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(data_in[15]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(data_in[1]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(data_in[2]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 output36 (.A(net36),
    .X(data_R));
 sky130_fd_sc_hd__buf_1 output37 (.A(net37),
    .X(data_W));
 sky130_fd_sc_hd__buf_1 output38 (.A(net38),
    .X(data_address[0]));
 sky130_fd_sc_hd__buf_1 output39 (.A(net39),
    .X(data_address[1]));
 sky130_fd_sc_hd__buf_1 output40 (.A(net40),
    .X(data_address[2]));
 sky130_fd_sc_hd__buf_1 output41 (.A(net41),
    .X(data_address[3]));
 sky130_fd_sc_hd__buf_1 output42 (.A(net42),
    .X(data_address[4]));
 sky130_fd_sc_hd__buf_1 output43 (.A(net43),
    .X(data_address[5]));
 sky130_fd_sc_hd__buf_1 output44 (.A(net44),
    .X(data_address[6]));
 sky130_fd_sc_hd__buf_1 output45 (.A(net45),
    .X(data_address[7]));
 sky130_fd_sc_hd__buf_1 output46 (.A(net46),
    .X(data_address[8]));
 sky130_fd_sc_hd__buf_1 output47 (.A(net47),
    .X(data_address[9]));
 sky130_fd_sc_hd__buf_1 output48 (.A(net48),
    .X(data_out[0]));
 sky130_fd_sc_hd__buf_1 output49 (.A(net49),
    .X(data_out[10]));
 sky130_fd_sc_hd__buf_1 output50 (.A(net50),
    .X(data_out[11]));
 sky130_fd_sc_hd__buf_1 output51 (.A(net51),
    .X(data_out[12]));
 sky130_fd_sc_hd__buf_1 output52 (.A(net52),
    .X(data_out[13]));
 sky130_fd_sc_hd__buf_1 output53 (.A(net53),
    .X(data_out[14]));
 sky130_fd_sc_hd__buf_1 output54 (.A(net54),
    .X(data_out[15]));
 sky130_fd_sc_hd__buf_1 output55 (.A(net55),
    .X(data_out[1]));
 sky130_fd_sc_hd__buf_1 output56 (.A(net56),
    .X(data_out[2]));
 sky130_fd_sc_hd__buf_1 output57 (.A(net57),
    .X(data_out[3]));
 sky130_fd_sc_hd__buf_1 output58 (.A(net58),
    .X(data_out[4]));
 sky130_fd_sc_hd__buf_1 output59 (.A(net59),
    .X(data_out[5]));
 sky130_fd_sc_hd__buf_1 output60 (.A(net60),
    .X(data_out[6]));
 sky130_fd_sc_hd__buf_1 output61 (.A(net61),
    .X(data_out[7]));
 sky130_fd_sc_hd__buf_1 output62 (.A(net62),
    .X(data_out[8]));
 sky130_fd_sc_hd__buf_1 output63 (.A(net63),
    .X(data_out[9]));
 sky130_fd_sc_hd__buf_1 output64 (.A(net64),
    .X(done));
 sky130_fd_sc_hd__buf_1 output65 (.A(net65),
    .X(instruction_address[0]));
 sky130_fd_sc_hd__buf_1 output66 (.A(net66),
    .X(instruction_address[1]));
 sky130_fd_sc_hd__buf_1 output67 (.A(net67),
    .X(instruction_address[2]));
 sky130_fd_sc_hd__buf_1 output68 (.A(net68),
    .X(instruction_address[3]));
 sky130_fd_sc_hd__buf_1 output69 (.A(net69),
    .X(instruction_address[4]));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net70),
    .X(instruction_address[5]));
 sky130_fd_sc_hd__buf_1 output71 (.A(net71),
    .X(instruction_address[6]));
 sky130_fd_sc_hd__buf_1 output72 (.A(net72),
    .X(instruction_address[7]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net73),
    .X(instruction_address[8]));
 sky130_fd_sc_hd__buf_1 output74 (.A(net74),
    .X(instruction_address[9]));
endmodule

