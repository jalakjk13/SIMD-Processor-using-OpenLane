VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO simd
  CLASS BLOCK ;
  FOREIGN simd ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 12.760 5.200 14.760 294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 42.760 5.200 44.760 294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 72.760 5.200 74.760 294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 102.760 5.200 104.760 294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 132.760 5.200 134.760 294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 162.760 5.200 164.760 294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 192.760 5.200 194.760 294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 222.760 5.200 224.760 294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 252.760 5.200 254.760 294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 282.760 5.200 284.760 294.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 13.140 295.100 15.140 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 43.140 295.100 45.140 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 73.140 295.100 75.140 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 103.140 295.100 105.140 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 133.140 295.100 135.140 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 163.140 295.100 165.140 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 193.140 295.100 195.140 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 223.140 295.100 225.140 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 253.140 295.100 255.140 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 283.140 295.100 285.140 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.060 5.200 11.060 294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.060 5.200 41.060 294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.060 5.200 71.060 294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.060 5.200 101.060 294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 129.060 5.200 131.060 294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 159.060 5.200 161.060 294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 189.060 5.200 191.060 294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 219.060 5.200 221.060 294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 249.060 5.200 251.060 294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 279.060 5.200 281.060 294.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 9.440 295.100 11.440 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 39.440 295.100 41.440 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 69.440 295.100 71.440 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 99.440 295.100 101.440 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 129.440 295.100 131.440 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 159.440 295.100 161.440 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 189.440 295.100 191.440 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 219.440 295.100 221.440 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 249.440 295.100 251.440 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 279.440 295.100 281.440 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 24.010 296.000 24.290 300.000 ;
    END
  END clk
  PIN data_R
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END data_R
  PIN data_W
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END data_W
  PIN data_address[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 156.440 300.000 157.040 ;
    END
  END data_address[0]
  PIN data_address[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 171.400 300.000 172.000 ;
    END
  END data_address[1]
  PIN data_address[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 186.360 300.000 186.960 ;
    END
  END data_address[2]
  PIN data_address[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 201.320 300.000 201.920 ;
    END
  END data_address[3]
  PIN data_address[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 216.280 300.000 216.880 ;
    END
  END data_address[4]
  PIN data_address[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 231.240 300.000 231.840 ;
    END
  END data_address[5]
  PIN data_address[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 246.200 300.000 246.800 ;
    END
  END data_address[6]
  PIN data_address[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 261.160 300.000 261.760 ;
    END
  END data_address[7]
  PIN data_address[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 276.120 300.000 276.720 ;
    END
  END data_address[8]
  PIN data_address[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 291.080 300.000 291.680 ;
    END
  END data_address[9]
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 55.290 296.000 55.570 300.000 ;
    END
  END data_in[0]
  PIN data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 211.690 296.000 211.970 300.000 ;
    END
  END data_in[10]
  PIN data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 227.330 296.000 227.610 300.000 ;
    END
  END data_in[11]
  PIN data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 242.970 296.000 243.250 300.000 ;
    END
  END data_in[12]
  PIN data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 258.610 296.000 258.890 300.000 ;
    END
  END data_in[13]
  PIN data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 274.250 296.000 274.530 300.000 ;
    END
  END data_in[14]
  PIN data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 289.890 296.000 290.170 300.000 ;
    END
  END data_in[15]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 70.930 296.000 71.210 300.000 ;
    END
  END data_in[1]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 86.570 296.000 86.850 300.000 ;
    END
  END data_in[2]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 102.210 296.000 102.490 300.000 ;
    END
  END data_in[3]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 117.850 296.000 118.130 300.000 ;
    END
  END data_in[4]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 133.490 296.000 133.770 300.000 ;
    END
  END data_in[5]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 149.130 296.000 149.410 300.000 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 164.770 296.000 165.050 300.000 ;
    END
  END data_in[7]
  PIN data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 180.410 296.000 180.690 300.000 ;
    END
  END data_in[8]
  PIN data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 196.050 296.000 196.330 300.000 ;
    END
  END data_in[9]
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END data_out[0]
  PIN data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END data_out[10]
  PIN data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END data_out[11]
  PIN data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END data_out[12]
  PIN data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END data_out[13]
  PIN data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END data_out[14]
  PIN data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END data_out[15]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END data_out[1]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END data_out[2]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END data_out[7]
  PIN data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END data_out[8]
  PIN data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END data_out[9]
  PIN done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END done
  PIN instruction_address[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 6.840 300.000 7.440 ;
    END
  END instruction_address[0]
  PIN instruction_address[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 21.800 300.000 22.400 ;
    END
  END instruction_address[1]
  PIN instruction_address[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 36.760 300.000 37.360 ;
    END
  END instruction_address[2]
  PIN instruction_address[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 51.720 300.000 52.320 ;
    END
  END instruction_address[3]
  PIN instruction_address[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 66.680 300.000 67.280 ;
    END
  END instruction_address[4]
  PIN instruction_address[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 81.640 300.000 82.240 ;
    END
  END instruction_address[5]
  PIN instruction_address[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 96.600 300.000 97.200 ;
    END
  END instruction_address[6]
  PIN instruction_address[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 111.560 300.000 112.160 ;
    END
  END instruction_address[7]
  PIN instruction_address[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 126.520 300.000 127.120 ;
    END
  END instruction_address[8]
  PIN instruction_address[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 296.000 141.480 300.000 142.080 ;
    END
  END instruction_address[9]
  PIN instruction_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END instruction_in[0]
  PIN instruction_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END instruction_in[10]
  PIN instruction_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END instruction_in[11]
  PIN instruction_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END instruction_in[12]
  PIN instruction_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END instruction_in[13]
  PIN instruction_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END instruction_in[14]
  PIN instruction_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END instruction_in[15]
  PIN instruction_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END instruction_in[16]
  PIN instruction_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END instruction_in[17]
  PIN instruction_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END instruction_in[1]
  PIN instruction_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END instruction_in[2]
  PIN instruction_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END instruction_in[3]
  PIN instruction_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END instruction_in[4]
  PIN instruction_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END instruction_in[5]
  PIN instruction_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END instruction_in[6]
  PIN instruction_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END instruction_in[7]
  PIN instruction_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END instruction_in[8]
  PIN instruction_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END instruction_in[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 39.650 296.000 39.930 300.000 ;
    END
  END rst
  OBS
      LAYER li1 ;
        RECT 5.060 5.355 294.860 293.845 ;
      LAYER met1 ;
        RECT 4.670 4.460 296.630 295.760 ;
      LAYER met2 ;
        RECT 4.690 295.720 23.730 296.210 ;
        RECT 24.570 295.720 39.370 296.210 ;
        RECT 40.210 295.720 55.010 296.210 ;
        RECT 55.850 295.720 70.650 296.210 ;
        RECT 71.490 295.720 86.290 296.210 ;
        RECT 87.130 295.720 101.930 296.210 ;
        RECT 102.770 295.720 117.570 296.210 ;
        RECT 118.410 295.720 133.210 296.210 ;
        RECT 134.050 295.720 148.850 296.210 ;
        RECT 149.690 295.720 164.490 296.210 ;
        RECT 165.330 295.720 180.130 296.210 ;
        RECT 180.970 295.720 195.770 296.210 ;
        RECT 196.610 295.720 211.410 296.210 ;
        RECT 212.250 295.720 227.050 296.210 ;
        RECT 227.890 295.720 242.690 296.210 ;
        RECT 243.530 295.720 258.330 296.210 ;
        RECT 259.170 295.720 273.970 296.210 ;
        RECT 274.810 295.720 289.610 296.210 ;
        RECT 290.450 295.720 296.600 296.210 ;
        RECT 4.690 4.280 296.600 295.720 ;
        RECT 4.690 3.670 23.730 4.280 ;
        RECT 24.570 3.670 38.450 4.280 ;
        RECT 39.290 3.670 53.170 4.280 ;
        RECT 54.010 3.670 67.890 4.280 ;
        RECT 68.730 3.670 82.610 4.280 ;
        RECT 83.450 3.670 97.330 4.280 ;
        RECT 98.170 3.670 112.050 4.280 ;
        RECT 112.890 3.670 126.770 4.280 ;
        RECT 127.610 3.670 141.490 4.280 ;
        RECT 142.330 3.670 156.210 4.280 ;
        RECT 157.050 3.670 170.930 4.280 ;
        RECT 171.770 3.670 185.650 4.280 ;
        RECT 186.490 3.670 200.370 4.280 ;
        RECT 201.210 3.670 215.090 4.280 ;
        RECT 215.930 3.670 229.810 4.280 ;
        RECT 230.650 3.670 244.530 4.280 ;
        RECT 245.370 3.670 259.250 4.280 ;
        RECT 260.090 3.670 273.970 4.280 ;
        RECT 274.810 3.670 288.690 4.280 ;
        RECT 289.530 3.670 296.600 4.280 ;
      LAYER met3 ;
        RECT 3.990 292.080 296.175 293.925 ;
        RECT 3.990 290.680 295.600 292.080 ;
        RECT 3.990 285.280 296.175 290.680 ;
        RECT 4.400 283.880 296.175 285.280 ;
        RECT 3.990 277.120 296.175 283.880 ;
        RECT 3.990 275.720 295.600 277.120 ;
        RECT 3.990 270.320 296.175 275.720 ;
        RECT 4.400 268.920 296.175 270.320 ;
        RECT 3.990 262.160 296.175 268.920 ;
        RECT 3.990 260.760 295.600 262.160 ;
        RECT 3.990 255.360 296.175 260.760 ;
        RECT 4.400 253.960 296.175 255.360 ;
        RECT 3.990 247.200 296.175 253.960 ;
        RECT 3.990 245.800 295.600 247.200 ;
        RECT 3.990 240.400 296.175 245.800 ;
        RECT 4.400 239.000 296.175 240.400 ;
        RECT 3.990 232.240 296.175 239.000 ;
        RECT 3.990 230.840 295.600 232.240 ;
        RECT 3.990 225.440 296.175 230.840 ;
        RECT 4.400 224.040 296.175 225.440 ;
        RECT 3.990 217.280 296.175 224.040 ;
        RECT 3.990 215.880 295.600 217.280 ;
        RECT 3.990 210.480 296.175 215.880 ;
        RECT 4.400 209.080 296.175 210.480 ;
        RECT 3.990 202.320 296.175 209.080 ;
        RECT 3.990 200.920 295.600 202.320 ;
        RECT 3.990 195.520 296.175 200.920 ;
        RECT 4.400 194.120 296.175 195.520 ;
        RECT 3.990 187.360 296.175 194.120 ;
        RECT 3.990 185.960 295.600 187.360 ;
        RECT 3.990 180.560 296.175 185.960 ;
        RECT 4.400 179.160 296.175 180.560 ;
        RECT 3.990 172.400 296.175 179.160 ;
        RECT 3.990 171.000 295.600 172.400 ;
        RECT 3.990 165.600 296.175 171.000 ;
        RECT 4.400 164.200 296.175 165.600 ;
        RECT 3.990 157.440 296.175 164.200 ;
        RECT 3.990 156.040 295.600 157.440 ;
        RECT 3.990 150.640 296.175 156.040 ;
        RECT 4.400 149.240 296.175 150.640 ;
        RECT 3.990 142.480 296.175 149.240 ;
        RECT 3.990 141.080 295.600 142.480 ;
        RECT 3.990 135.680 296.175 141.080 ;
        RECT 4.400 134.280 296.175 135.680 ;
        RECT 3.990 127.520 296.175 134.280 ;
        RECT 3.990 126.120 295.600 127.520 ;
        RECT 3.990 120.720 296.175 126.120 ;
        RECT 4.400 119.320 296.175 120.720 ;
        RECT 3.990 112.560 296.175 119.320 ;
        RECT 3.990 111.160 295.600 112.560 ;
        RECT 3.990 105.760 296.175 111.160 ;
        RECT 4.400 104.360 296.175 105.760 ;
        RECT 3.990 97.600 296.175 104.360 ;
        RECT 3.990 96.200 295.600 97.600 ;
        RECT 3.990 90.800 296.175 96.200 ;
        RECT 4.400 89.400 296.175 90.800 ;
        RECT 3.990 82.640 296.175 89.400 ;
        RECT 3.990 81.240 295.600 82.640 ;
        RECT 3.990 75.840 296.175 81.240 ;
        RECT 4.400 74.440 296.175 75.840 ;
        RECT 3.990 67.680 296.175 74.440 ;
        RECT 3.990 66.280 295.600 67.680 ;
        RECT 3.990 60.880 296.175 66.280 ;
        RECT 4.400 59.480 296.175 60.880 ;
        RECT 3.990 52.720 296.175 59.480 ;
        RECT 3.990 51.320 295.600 52.720 ;
        RECT 3.990 45.920 296.175 51.320 ;
        RECT 4.400 44.520 296.175 45.920 ;
        RECT 3.990 37.760 296.175 44.520 ;
        RECT 3.990 36.360 295.600 37.760 ;
        RECT 3.990 30.960 296.175 36.360 ;
        RECT 4.400 29.560 296.175 30.960 ;
        RECT 3.990 22.800 296.175 29.560 ;
        RECT 3.990 21.400 295.600 22.800 ;
        RECT 3.990 7.840 296.175 21.400 ;
        RECT 3.990 6.440 295.600 7.840 ;
        RECT 3.990 4.935 296.175 6.440 ;
      LAYER met4 ;
        RECT 17.775 4.935 38.660 292.905 ;
        RECT 41.460 4.935 42.360 292.905 ;
        RECT 45.160 4.935 68.660 292.905 ;
        RECT 71.460 4.935 72.360 292.905 ;
        RECT 75.160 4.935 98.660 292.905 ;
        RECT 101.460 4.935 102.360 292.905 ;
        RECT 105.160 4.935 128.660 292.905 ;
        RECT 131.460 4.935 132.360 292.905 ;
        RECT 135.160 4.935 158.660 292.905 ;
        RECT 161.460 4.935 162.360 292.905 ;
        RECT 165.160 4.935 188.660 292.905 ;
        RECT 191.460 4.935 192.360 292.905 ;
        RECT 195.160 4.935 218.660 292.905 ;
        RECT 221.460 4.935 222.360 292.905 ;
        RECT 225.160 4.935 248.660 292.905 ;
        RECT 251.460 4.935 252.360 292.905 ;
        RECT 255.160 4.935 278.660 292.905 ;
        RECT 281.460 4.935 282.360 292.905 ;
        RECT 285.160 4.935 291.345 292.905 ;
      LAYER met5 ;
        RECT 18.980 256.740 289.220 274.500 ;
        RECT 18.980 226.740 289.220 247.840 ;
        RECT 18.980 196.740 289.220 217.840 ;
        RECT 18.980 166.740 289.220 187.840 ;
        RECT 18.980 136.740 289.220 157.840 ;
        RECT 18.980 106.740 289.220 127.840 ;
        RECT 18.980 79.100 289.220 97.840 ;
  END
END simd
END LIBRARY

