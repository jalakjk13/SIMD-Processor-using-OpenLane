* NGSPICE file created from simd.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

.subckt simd VGND VPWR clk data_R data_W data_address[0] data_address[1] data_address[2]
+ data_address[3] data_address[4] data_address[5] data_address[6] data_address[7]
+ data_address[8] data_address[9] data_in[0] data_in[10] data_in[11] data_in[12] data_in[13]
+ data_in[14] data_in[15] data_in[1] data_in[2] data_in[3] data_in[4] data_in[5] data_in[6]
+ data_in[7] data_in[8] data_in[9] data_out[0] data_out[10] data_out[11] data_out[12]
+ data_out[13] data_out[14] data_out[15] data_out[1] data_out[2] data_out[3] data_out[4]
+ data_out[5] data_out[6] data_out[7] data_out[8] data_out[9] done instruction_address[0]
+ instruction_address[1] instruction_address[2] instruction_address[3] instruction_address[4]
+ instruction_address[5] instruction_address[6] instruction_address[7] instruction_address[8]
+ instruction_address[9] instruction_in[0] instruction_in[10] instruction_in[11] instruction_in[12]
+ instruction_in[13] instruction_in[14] instruction_in[15] instruction_in[16] instruction_in[17]
+ instruction_in[1] instruction_in[2] instruction_in[3] instruction_in[4] instruction_in[5]
+ instruction_in[6] instruction_in[7] instruction_in[8] instruction_in[9] rst
XFILLER_0_94_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06883_ result_reg_mac\[12\] VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__inv_2
X_09671_ Oset\[3\]\[6\] _03024_ _03026_ VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08622_ _02532_ _02535_ _02536_ VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__nand3_1
X_08553_ _02470_ H\[0\]\[13\] VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07504_ _01568_ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08484_ _02404_ net49 _02169_ VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07435_ result_reg_mac\[14\] _01215_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07366_ result_reg_not\[11\] _01439_ _01167_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07297_ _00881_ _01374_ _01182_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06317_ LC\[5\] _06277_ VGND VGND VPWR VPWR _06278_ sky130_fd_sc_hd__nor2_1
X_09105_ _02556_ _03015_ VGND VGND VPWR VPWR _03016_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09036_ _02947_ _02237_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09938_ _03157_ Oset\[3\]\[9\] _03135_ _03844_ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__a211o_1
XFILLER_0_99_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09869_ Qset\[3\]\[8\] _03341_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__nor2_1
X_12880_ clknet_leaf_20_clk _00323_ VGND VGND VPWR VPWR result_reg_Lshift\[15\] sky130_fd_sc_hd__dfxtp_1
X_11900_ _02790_ _02793_ VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__nand2_2
XFILLER_0_68_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11831_ _05699_ VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11762_ _05627_ _04642_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11693_ _05554_ _04830_ _05592_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__nand3_1
X_10713_ Qset\[1\]\[10\] _03791_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__nand2_1
X_10644_ _04105_ Qset\[3\]\[10\] _04045_ _04548_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_11_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10575_ _04282_ Oset\[2\]\[10\] _03345_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__o21ai_1
X_12314_ _06055_ _00930_ VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12245_ _06031_ VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__clkbuf_4
X_12176_ _05974_ _00524_ _05937_ _05975_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__a22o_1
X_11127_ _05014_ _05012_ _05013_ _04954_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__o2bb2a_1
X_11058_ _04881_ _02455_ VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__nor2_1
X_10009_ _03912_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07220_ _00770_ _01267_ _01263_ _01301_ VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__a211o_1
XFILLER_0_73_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07151_ _00528_ _00631_ _00634_ _01171_ VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__or4_1
XFILLER_0_54_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07082_ _01163_ _00654_ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_74_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07984_ _02004_ VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__clkbuf_1
X_06935_ result_reg_mac\[14\] VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__inv_2
X_09723_ _03498_ Oset\[1\]\[7\] _02991_ _03630_ VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__a211o_1
X_06866_ _00989_ _00553_ VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__or2_1
X_09654_ _03560_ _03537_ _03540_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__nand3_1
X_08605_ _02520_ net54 _02169_ VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__mux2_1
X_06797_ _00922_ _00923_ _00643_ VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__mux2_1
X_09585_ _02302_ _00584_ VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__nand2_1
X_08536_ _02397_ Qset\[3\]\[13\] _02374_ _02453_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08467_ _02356_ _02387_ VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__nor2_1
X_07418_ _01276_ _01476_ _01488_ _01489_ VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__a22o_2
X_08398_ _02319_ Oset\[3\]\[7\] _02254_ _02321_ VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__a211o_1
X_07349_ net2 _01255_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10360_ _04204_ _04265_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__nor2_1
X_10291_ _04195_ _04196_ _04197_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__nand3_2
X_09019_ _02586_ Qset\[1\]\[3\] VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__nand2_1
X_12030_ result_reg_Rshift\[6\] _05848_ _05857_ _05858_ VGND VGND VPWR VPWR _00330_
+ sky130_fd_sc_hd__o211a_1
X_12932_ clknet_leaf_22_clk _00375_ VGND VGND VPWR VPWR result_reg_not\[3\] sky130_fd_sc_hd__dfxtp_1
X_12863_ clknet_leaf_10_clk _00306_ VGND VGND VPWR VPWR result_reg_mac\[14\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_44_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11814_ _05688_ VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__inv_2
X_12794_ clknet_leaf_44_clk _00237_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dfxtp_1
X_11745_ _00788_ _05631_ _05634_ _05639_ VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11676_ _05517_ _02577_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_24_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10627_ _04040_ _04365_ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_11_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10558_ _04459_ _04462_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__or2_1
X_12228_ _05141_ _04969_ _05881_ VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__a21o_1
X_10489_ _04391_ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12159_ _05960_ _05961_ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06720_ result_reg_Lshift\[5\] VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__inv_2
X_06651_ _00777_ _00782_ VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__nand2_4
XFILLER_0_91_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06582_ _00702_ _00703_ _00539_ VGND VGND VPWR VPWR _00716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09370_ _03280_ Add.sub VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08321_ _02141_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__buf_4
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08252_ Oset\[0\]\[1\] VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07203_ _01282_ _01207_ _01261_ _01285_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08183_ _02115_ VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__buf_4
XFILLER_0_61_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07134_ _00661_ _00654_ _01163_ VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_42_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07065_ R0\[1\] net19 current_state\[2\] VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07967_ _01960_ _06281_ _01986_ VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__o21a_1
X_06918_ _01032_ _00600_ _01039_ _00699_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09706_ _03613_ VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__inv_2
X_07898_ Oset\[2\]\[2\] _01295_ _01942_ VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06849_ result_reg_not\[10\] VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09637_ _03110_ _03020_ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__nand2_1
X_09568_ _03475_ _03476_ VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08519_ _02364_ Oset\[3\]\[12\] _02347_ _02437_ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__a211o_1
X_11530_ _05412_ _05430_ VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__nand2_1
X_09499_ _03406_ VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11461_ _05065_ _05236_ _05240_ VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_21_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11392_ _05292_ _05293_ VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__nand2_1
X_10412_ _04262_ _04317_ VGND VGND VPWR VPWR _04318_ sky130_fd_sc_hd__nand2_2
X_10343_ _00710_ _03835_ _04249_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_94_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10274_ _04163_ _04178_ _04180_ VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__o21ai_1
X_12013_ _05843_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12915_ clknet_leaf_15_clk _00358_ VGND VGND VPWR VPWR result_reg_or\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_57_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12846_ clknet_leaf_4_clk _00289_ VGND VGND VPWR VPWR result_reg_mul\[13\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12777_ clknet_leaf_25_clk _00220_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11728_ _05626_ VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11659_ _05362_ _05368_ _05372_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08870_ _02776_ _02782_ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__nand2_1
X_07821_ _01594_ _01866_ _01873_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__o21ai_1
X_07752_ _00939_ _01574_ _01569_ _01807_ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__a211o_1
X_07683_ _00865_ _00857_ _01545_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__mux2_1
X_06703_ CMD_addition VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__inv_2
X_06634_ _00765_ _00745_ VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__or2_1
X_09422_ _03001_ Oset\[3\]\[5\] VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09353_ _03237_ _03263_ VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__nor2_1
X_06565_ _00697_ _00605_ _00698_ _00606_ VGND VGND VPWR VPWR _00699_ sky130_fd_sc_hd__or4_4
X_08304_ H\[3\]\[3\] _02230_ VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06496_ current_state\[5\] VGND VGND VPWR VPWR _00631_ sky130_fd_sc_hd__buf_2
X_09284_ _03191_ _03193_ _03194_ VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08235_ _02165_ _02123_ VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08166_ _02102_ _02103_ net40 VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__a21o_1
X_07117_ _01201_ VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__buf_4
X_08097_ _01781_ H\[1\]\[7\] _02057_ VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07048_ _01140_ VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08999_ _02736_ _02823_ VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10961_ _02446_ _04856_ _04863_ VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12700_ clknet_leaf_26_clk _00150_ VGND VGND VPWR VPWR Oset\[0\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10892_ _04792_ _00831_ _04793_ VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__nand3_1
X_12631_ clknet_leaf_41_clk _00081_ VGND VGND VPWR VPWR Oset\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12562_ _06085_ _05134_ VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11513_ _05209_ _05212_ _05211_ VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__a21oi_1
X_12493_ _06212_ VGND VGND VPWR VPWR _00439_ sky130_fd_sc_hd__clkbuf_1
X_11444_ _02494_ _04856_ _05344_ VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11375_ _05275_ _05276_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__nand2_1
X_10326_ _04222_ _04232_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10257_ _03920_ _03956_ _03919_ VGND VGND VPWR VPWR _04164_ sky130_fd_sc_hd__a21oi_1
X_10188_ _04088_ _04094_ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_6_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12829_ clknet_leaf_9_clk _00272_ VGND VGND VPWR VPWR result_reg_sub\[12\] sky130_fd_sc_hd__dfxtp_1
X_06350_ _00484_ _00490_ VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_60_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08020_ _02023_ VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09971_ _03869_ _03877_ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__or2_1
X_08922_ _02833_ _02834_ VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__nand2_1
X_08853_ _02764_ _00005_ _02765_ VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__nand3_1
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07804_ result_reg_not\[11\] _01633_ _01857_ VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__a21o_1
X_08784_ Oset\[3\]\[1\] _02625_ _02626_ _02697_ VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__a211o_1
X_07735_ _01789_ _01663_ _01790_ _01791_ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_68_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07666_ net12 _01658_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__nor2_1
X_09405_ _02822_ _03308_ VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__nor2_1
X_06617_ _00737_ _00619_ _00629_ _00749_ VGND VGND VPWR VPWR _00750_ sky130_fd_sc_hd__a211o_1
X_07597_ _01655_ _01635_ _01657_ _01659_ VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__a31o_1
XFILLER_0_94_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06548_ _00498_ _00629_ _00680_ _00682_ _00664_ VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__a221o_1
X_09336_ _03243_ VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09267_ _03177_ VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06479_ _00609_ _00612_ _00613_ VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__mux2_1
X_08218_ _02131_ _02146_ _02147_ _02148_ VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_15_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09198_ _03078_ _03108_ VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__nand2_1
X_08149_ Add.sub VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_91_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11160_ _03790_ _03745_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__nand2_1
X_11091_ _04975_ _04691_ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__nor2_1
X_10111_ _04016_ _04017_ VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10042_ _03897_ _03899_ _02620_ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__or3b_1
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11993_ _05831_ VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10944_ _04843_ _04844_ _04845_ _04846_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__o22a_1
X_10875_ _04778_ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12614_ clknet_leaf_40_clk _00064_ VGND VGND VPWR VPWR Qset\[2\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12545_ _06243_ VGND VGND VPWR VPWR _00460_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12476_ _06199_ _01146_ _06201_ VGND VGND VPWR VPWR _06202_ sky130_fd_sc_hd__and3_1
XANTENNA_5 _00567_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11427_ _05319_ Qset\[1\]\[14\] _04835_ _05327_ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__a211o_1
X_11358_ _04690_ _04460_ VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10309_ _03897_ _02578_ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__nor2_1
X_11289_ _05188_ _05187_ VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07520_ _01584_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_65_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07451_ _01520_ _01187_ VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06402_ _00536_ CMD_addition _06264_ _00529_ VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__or4_4
X_07382_ Oset\[3\]\[11\] _01455_ _01249_ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06333_ _00477_ VGND VGND VPWR VPWR _00478_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09121_ _03022_ Qset\[0\]\[4\] VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09052_ _02836_ _02231_ VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08003_ Oset\[0\]\[12\] _01473_ _02000_ VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09954_ H\[0\]\[11\] VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__inv_2
X_08905_ _02817_ _02572_ _00586_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__a21oi_1
X_09885_ _03791_ VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08836_ _02748_ _02749_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__and2_2
X_08767_ _02678_ _02680_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07718_ result_reg_and\[7\] VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__inv_2
X_08698_ _02611_ H\[3\]\[0\] _02591_ _02612_ VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__a211o_1
X_07649_ result_reg_mul\[4\] _01688_ _01589_ VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10660_ _04563_ _04537_ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09319_ _03214_ _03216_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10591_ _04281_ _04495_ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12330_ R3\[1\] net26 current_state\[2\] VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12261_ _06039_ _05785_ _06013_ _06041_ VGND VGND VPWR VPWR _00378_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11212_ _05113_ _03746_ _05114_ VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__nand3_2
Xoutput42 net42 VGND VGND VPWR VPWR data_address[4] sky130_fd_sc_hd__buf_1
X_12192_ _05783_ _03489_ _05907_ VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11143_ _04992_ _05045_ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__nand2_1
Xoutput64 net64 VGND VGND VPWR VPWR done sky130_fd_sc_hd__buf_1
Xoutput53 net53 VGND VGND VPWR VPWR data_out[14] sky130_fd_sc_hd__buf_1
XFILLER_0_37_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11074_ _04959_ _04976_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__nand2b_1
X_10025_ _03929_ _03931_ VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _00590_ _04741_ _04735_ _01158_ _05816_ VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__a221o_2
X_10927_ _00820_ VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__buf_6
XFILLER_0_73_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10858_ _04584_ _04575_ _04583_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_70_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10789_ _04667_ _04692_ VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_14_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12528_ _00668_ Qset\[3\]\[0\] _06234_ VGND VGND VPWR VPWR _06235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12459_ _06188_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06951_ net6 _00735_ _00839_ _01071_ VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__o211a_1
X_09670_ Oset\[1\]\[6\] _03024_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06882_ _01005_ VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__clkbuf_1
X_08621_ Qset\[1\]\[0\] _02529_ VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08552_ _02459_ VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__buf_4
X_07503_ _01567_ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08483_ _02139_ _02390_ _02126_ _02395_ _02403_ VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__o221ai_4
X_07434_ _01503_ _01261_ _01190_ _01504_ VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__a211o_1
X_07365_ result_reg_Lshift\[11\] result_reg_Rshift\[11\] _01164_ VGND VGND VPWR VPWR
+ _01439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07296_ _00882_ _01373_ _01177_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06316_ _06276_ VGND VGND VPWR VPWR _06277_ sky130_fd_sc_hd__inv_2
X_09104_ _03011_ _03012_ _03013_ _03014_ VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__o22a_1
XFILLER_0_32_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09035_ _02946_ _01552_ VGND VGND VPWR VPWR _02947_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09937_ _02545_ _02365_ VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__nor2_1
X_09868_ _03345_ _03771_ _03772_ _03774_ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_99_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09799_ _03705_ _03706_ VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__nand2_1
X_08819_ _00586_ R3\[1\] VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__nand2_1
X_11830_ _05673_ _05470_ _05698_ VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__o21ai_1
X_11761_ _05650_ VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__inv_2
Xclkbuf_3_6__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10712_ _03023_ Qset\[0\]\[10\] VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__nand2_1
X_11692_ _05555_ _05590_ _05591_ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_36_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10643_ _04105_ _04472_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10574_ Oset\[3\]\[10\] _03773_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12313_ _05766_ _00669_ _03857_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12244_ _06030_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_31_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12175_ _02881_ _02923_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__nand2_1
X_11126_ _04495_ _04899_ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__nor2_1
X_11057_ Qset\[2\]\[13\] Qset\[3\]\[13\] _04729_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10008_ _03886_ _03891_ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_47_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11959_ _05774_ _05801_ _05672_ _05802_ VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__o211a_1
X_07150_ _00557_ current_state\[5\] _00634_ _01234_ VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__or4_1
XFILLER_0_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07081_ result_reg_Lshift\[0\] result_reg_Rshift\[0\] _01165_ VGND VGND VPWR VPWR
+ _01166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07983_ Oset\[0\]\[2\] _01295_ _02001_ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__mux2_1
X_09722_ _03498_ _02323_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__nor2_1
X_06934_ _01055_ VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06865_ result_reg_or\[11\] VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__inv_2
X_09653_ _03541_ _03561_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__nand2_1
X_08604_ _02311_ _02506_ _02139_ _02513_ _02519_ VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__o221ai_4
X_09584_ _03484_ _03492_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__nand2_1
X_06796_ result_reg_Lshift\[8\] VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__inv_2
X_08535_ _02397_ _02452_ VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08466_ Oset\[0\]\[10\] VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__inv_2
X_07417_ _01031_ _01275_ _01160_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__a21oi_1
X_08397_ _02261_ _02320_ VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__nor2_1
X_07348_ result_reg_not\[10\] _01422_ _01167_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07279_ _01356_ _01193_ _01192_ _01357_ VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__a211o_1
XFILLER_0_60_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10290_ _04041_ _03751_ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__nand2_1
X_09018_ _02582_ Qset\[0\]\[3\] VGND VGND VPWR VPWR _02930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12931_ clknet_leaf_22_clk _00374_ VGND VGND VPWR VPWR result_reg_not\[2\] sky130_fd_sc_hd__dfxtp_1
X_12862_ clknet_leaf_9_clk _00305_ VGND VGND VPWR VPWR result_reg_mac\[13\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_87_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11813_ _04198_ _04248_ _05677_ _05687_ VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_44_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ clknet_leaf_44_clk _00236_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dfxtp_1
X_11744_ _05627_ _03293_ VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11675_ _05341_ _02734_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_99_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10626_ _04528_ _04530_ VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10557_ _04265_ _04461_ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10488_ _04040_ _04028_ _04363_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__nand3_1
X_12227_ result_reg_or\[12\] _05959_ _06013_ _06017_ VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__o211a_1
X_12158_ _02538_ _02595_ _05907_ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12089_ _01666_ VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__buf_4
X_11109_ _04975_ _04025_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__nor2_1
X_06650_ _00778_ _00655_ _00657_ _00781_ _00666_ VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06581_ result_reg_and\[1\] VGND VGND VPWR VPWR _00715_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08320_ _02243_ _02246_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08251_ _02131_ _02179_ _00003_ _02180_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_24_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07202_ _00727_ _01204_ _01245_ _01284_ VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08182_ _00635_ VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__buf_4
XFILLER_0_6_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07133_ _01161_ _01169_ _01217_ VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__a21bo_4
XFILLER_0_15_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07064_ _01150_ VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07966_ _01986_ _01991_ VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__nand2_1
X_06917_ _01033_ _01038_ _00607_ VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__mux2_1
X_09705_ _02895_ _03079_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__nand2_1
X_07897_ _01944_ VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__clkbuf_1
X_09636_ _03076_ _03020_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__nand2_1
X_06848_ _00955_ _00725_ _00972_ VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06779_ result_reg_add\[8\] VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__inv_2
X_09567_ _03473_ _03466_ _03470_ VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__nand3_1
XFILLER_0_65_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08518_ _02364_ _02436_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__nor2_1
X_09498_ _03231_ _03215_ _03214_ VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08449_ _02367_ _02370_ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__nand2_2
X_11460_ _05079_ _04495_ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_21_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11391_ _05291_ _05287_ _05288_ VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__nand3b_1
X_10411_ _04316_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10342_ _04198_ _04248_ _00710_ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__nand3_1
XFILLER_0_33_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12012_ _05844_ _05845_ _05808_ _05846_ VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__o211a_1
X_10273_ _04162_ _04179_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__or2_1
X_12914_ clknet_leaf_15_clk _00357_ VGND VGND VPWR VPWR result_reg_or\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_57_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12845_ clknet_leaf_4_clk _00288_ VGND VGND VPWR VPWR result_reg_mul\[12\] sky130_fd_sc_hd__dfxtp_1
X_12776_ clknet_leaf_27_clk _00219_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ CMD_addition _00832_ _06269_ VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__or3_1
XFILLER_0_56_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11658_ _05557_ _04190_ VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11589_ _05489_ VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10609_ _04454_ _04513_ VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_71_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07820_ _01870_ _01595_ _01871_ _01872_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__a31o_1
X_07751_ _01407_ _01577_ _01572_ _01806_ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__o211a_1
X_06702_ _00831_ VGND VGND VPWR VPWR _00832_ sky130_fd_sc_hd__buf_4
X_07682_ _01741_ VGND VGND VPWR VPWR _00099_ sky130_fd_sc_hd__clkbuf_1
X_06633_ result_reg_mul\[3\] VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__inv_2
X_09421_ _03329_ _03330_ _02540_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_82_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06564_ _00597_ _00578_ VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__nand2_1
X_09352_ _03260_ _03262_ VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__nand2_1
X_08303_ H\[2\]\[3\] VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__inv_2
X_06495_ _00564_ _00604_ _00618_ _00619_ _00629_ VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09283_ _03184_ _03145_ VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__nand2_1
X_08234_ _02160_ _02164_ VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__nor2_1
X_08165_ R3\[1\] _02100_ _02105_ _02106_ VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07116_ _01200_ _00537_ VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08096_ _02064_ VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07047_ _00979_ Qset\[2\]\[10\] _01128_ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08998_ _02902_ _02909_ VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__nand2_1
X_07949_ _06275_ LC\[4\] VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__and2_1
X_10960_ _04856_ H\[0\]\[12\] _04862_ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10891_ _04794_ _02160_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_26_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09619_ _03377_ _03376_ VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12630_ clknet_leaf_44_clk _00080_ VGND VGND VPWR VPWR Oset\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_12561_ _06251_ VGND VGND VPWR VPWR _00468_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11512_ _05218_ _05215_ VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__nand2_1
X_12492_ _01531_ _05134_ VGND VGND VPWR VPWR _06212_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11443_ _04856_ H\[0\]\[14\] _04862_ VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11374_ _05089_ _05102_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10325_ _04228_ _04231_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__nand2_1
X_10256_ _03986_ _04160_ _04162_ VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10187_ _04093_ _02573_ _00588_ VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_6_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12828_ clknet_leaf_10_clk _00271_ VGND VGND VPWR VPWR result_reg_sub\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12759_ clknet_leaf_49_clk _00202_ VGND VGND VPWR VPWR H\[0\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09970_ _02687_ _03876_ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__nand2_1
X_08921_ _02831_ _00536_ _02832_ VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__nand3_1
X_08852_ _02585_ Oset\[3\]\[2\] VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__nand2_1
X_07803_ result_reg_Rshift\[11\] _01672_ _01601_ _01856_ VGND VGND VPWR VPWR _01857_
+ sky130_fd_sc_hd__o211a_1
X_08783_ _02625_ _02179_ VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_49_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_8
X_07734_ result_reg_mul\[8\] _01688_ _01667_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_68_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07665_ _00840_ _01682_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__or2_1
X_06616_ _00738_ _00709_ _00739_ _00748_ VGND VGND VPWR VPWR _00749_ sky130_fd_sc_hd__o211a_1
X_09404_ _03310_ _03313_ VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__nand2_1
X_07596_ net9 _01658_ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__nor2_1
X_06547_ _00602_ _00681_ VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09335_ _02898_ _03245_ VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06478_ _00532_ _00574_ VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__nand2_4
XFILLER_0_62_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09266_ _03176_ _03116_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08217_ _02141_ Oset\[1\]\[0\] VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09197_ _03107_ VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__inv_2
X_08148_ _02091_ VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08079_ _02054_ VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11090_ _04992_ _04989_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__and2_1
X_10110_ _03652_ _03745_ _03859_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__nand3_1
X_10041_ _03947_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__inv_2
X_11992_ _05829_ _05771_ _05775_ _05830_ VGND VGND VPWR VPWR _05831_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_3_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10943_ Qset\[1\]\[12\] _03773_ _03004_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10874_ _04776_ _04777_ VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12613_ clknet_leaf_43_clk _00063_ VGND VGND VPWR VPWR Qset\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12544_ _00927_ Qset\[3\]\[8\] _06234_ VGND VGND VPWR VPWR _06243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12475_ _06130_ _06167_ _06106_ _06200_ VGND VGND VPWR VPWR _06201_ sky130_fd_sc_hd__o22a_1
X_11426_ _04832_ _02479_ VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_6 _00621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11357_ _04690_ _04651_ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10308_ _04213_ _04214_ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__nand2_1
X_11288_ _05189_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__inv_2
X_10239_ _04145_ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07450_ _01092_ _01519_ _01182_ VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__mux2_1
X_07381_ _01276_ _01440_ _01453_ _01454_ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__a22o_2
X_06401_ Add.sub VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06332_ _00473_ _06259_ VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__nand2_1
X_09120_ H\[0\]\[4\] _03023_ _03030_ VGND VGND VPWR VPWR _03031_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09051_ _02948_ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__buf_6
XFILLER_0_72_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08002_ _02013_ VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_77_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09953_ _03859_ _02963_ _03745_ VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__nand3_1
X_09884_ _03025_ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__clkbuf_4
X_08904_ _02813_ _02814_ _02816_ VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__o21ai_2
X_08835_ _02747_ _02744_ _02745_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__nand3_1
X_08766_ _02585_ H\[3\]\[1\] _02590_ _02679_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__a211o_1
X_07717_ _01772_ _01585_ _01773_ _01774_ VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_0_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ _02586_ _02152_ VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__nor2_1
X_07648_ _01586_ result_reg_sub\[4\] VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07579_ result_reg_mul\[1\] _01585_ _01589_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09318_ _03214_ _03216_ _03228_ VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10590_ _04494_ VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__inv_2
X_09249_ _02562_ Qset\[3\]\[4\] _02800_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12260_ _06033_ _00873_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__nand2_1
X_12191_ _05937_ _05986_ _05987_ _05904_ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__a22o_1
X_11211_ _05112_ _05055_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput43 net43 VGND VGND VPWR VPWR data_address[5] sky130_fd_sc_hd__buf_1
X_11142_ _04691_ _04899_ _04991_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_8_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput54 net54 VGND VGND VPWR VPWR data_out[15] sky130_fd_sc_hd__buf_1
Xoutput65 net65 VGND VGND VPWR VPWR instruction_address[0] sky130_fd_sc_hd__buf_1
X_11073_ _04958_ _04954_ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__nand2_1
X_10024_ _03930_ _03869_ VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_62_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11975_ _01554_ _03866_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10926_ _04829_ VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__inv_2
X_10857_ _04593_ _04589_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_70_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10788_ _04281_ _04691_ VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12527_ _06233_ VGND VGND VPWR VPWR _06234_ sky130_fd_sc_hd__clkbuf_8
X_12458_ _06164_ _06105_ VGND VGND VPWR VPWR _06188_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11409_ _05308_ _05310_ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__nor2_1
X_12389_ net20 VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06950_ _01070_ _00735_ VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06881_ _01004_ Qset\[0\]\[11\] _00686_ VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__mux2_1
X_08620_ _02534_ VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__clkbuf_8
X_08551_ H\[1\]\[13\] VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07502_ _01566_ _01559_ _01560_ VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08482_ _02399_ _02402_ _01553_ VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__a21o_2
X_07433_ result_reg_or\[14\] _01199_ VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07364_ _01438_ VGND VGND VPWR VPWR _00084_ sky130_fd_sc_hd__clkbuf_1
X_09103_ H\[1\]\[4\] _02582_ _02591_ VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__o21ai_1
X_07295_ _00883_ _00884_ _01174_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06315_ LC\[4\] _06275_ VGND VGND VPWR VPWR _06276_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09034_ _02938_ _02945_ VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09936_ _02565_ Oset\[1\]\[9\] _02526_ _03842_ VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__a211o_1
X_09867_ Oset\[1\]\[8\] _03773_ _03761_ VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09798_ _00623_ _03076_ VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__or2_1
X_08818_ _02724_ _02731_ VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08749_ _02178_ shift.Q VGND VGND VPWR VPWR _02663_ sky130_fd_sc_hd__nand2_1
X_11760_ _00932_ _05631_ _05634_ _05649_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10711_ _02400_ _04415_ _04615_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11691_ _05555_ _05590_ _04196_ VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__a21oi_1
X_10642_ _04546_ _03781_ _00585_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10573_ _04477_ _00582_ VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_11_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12312_ _06073_ _06055_ _06066_ _06074_ VGND VGND VPWR VPWR _00396_ sky130_fd_sc_hd__o211a_1
X_12243_ _02164_ _05955_ _02098_ _00632_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__or4_2
XPHY_EDGE_ROW_39_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12174_ _02933_ _05760_ VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__nand2_1
X_11125_ _05027_ _05024_ VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__nand2_1
X_11056_ _04954_ _04958_ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__nor2_1
X_10007_ _03913_ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_48_Left_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11958_ _05774_ _00901_ VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11889_ _05740_ VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10909_ _01538_ _04798_ _04800_ _00556_ _04812_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__a311o_2
X_07080_ _01164_ VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__buf_4
XFILLER_0_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07982_ _02003_ VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__clkbuf_1
X_06933_ _01054_ Qset\[0\]\[13\] _00686_ VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__mux2_1
X_09721_ _03498_ Oset\[3\]\[7\] _03004_ _03628_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__a211o_1
X_06864_ _00984_ _00743_ _00986_ _00987_ VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_66_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09652_ _03560_ VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06795_ result_reg_Rshift\[8\] VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__inv_2
X_08603_ _02516_ _02518_ _01554_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__a21o_1
X_09583_ _03490_ _03491_ _02540_ VGND VGND VPWR VPWR _03492_ sky130_fd_sc_hd__nand3_1
XFILLER_0_89_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08534_ Qset\[2\]\[13\] VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08465_ _02364_ Oset\[3\]\[10\] _02347_ _02385_ VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__a211o_1
X_07416_ _01254_ _01477_ _01481_ _01487_ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08396_ Oset\[2\]\[7\] VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__inv_2
X_07347_ result_reg_Lshift\[10\] result_reg_Rshift\[10\] _01164_ VGND VGND VPWR VPWR
+ _01422_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_75_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07278_ net13 _01193_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09017_ _02927_ _02584_ _02928_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__nand3_1
XFILLER_0_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_84_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09919_ _03820_ _03825_ _01155_ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__nand3_1
X_12930_ clknet_leaf_19_clk _00373_ VGND VGND VPWR VPWR result_reg_not\[1\] sky130_fd_sc_hd__dfxtp_1
X_12861_ clknet_leaf_8_clk _00304_ VGND VGND VPWR VPWR result_reg_mac\[12\] sky130_fd_sc_hd__dfxtp_2
X_11812_ result_reg_mul\[8\] _05669_ _05682_ VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_16_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ clknet_leaf_45_clk _00235_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dfxtp_1
X_11743_ _05638_ VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11674_ _05382_ _05385_ _05384_ VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_99_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10625_ _04529_ _04392_ _04396_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_91_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10556_ _03790_ _04460_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__nand2_1
X_10487_ _04340_ _04365_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__nand2_1
X_12226_ _05937_ _06014_ _06015_ _05957_ _06016_ VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__a2111o_1
X_12157_ _05958_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__buf_2
X_11108_ _04309_ _04899_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__nor2_1
X_12088_ _03003_ _03006_ VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__and2_1
X_11039_ _04940_ _04923_ VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06580_ _00713_ VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08250_ _02131_ Oset\[3\]\[1\] VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__nand2_1
X_07201_ _01204_ _01283_ VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__nor2_1
X_08181_ im_reg\[9\] _02100_ _02105_ _02114_ VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07132_ _01195_ _01212_ _01214_ _01160_ _01216_ VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__a311o_1
XFILLER_0_54_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07063_ _01147_ _01149_ VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07965_ _01960_ _01990_ _06280_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__a21o_1
X_06916_ _01034_ _01037_ _00613_ VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__mux2_1
X_09704_ _03421_ _03462_ VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07896_ Oset\[2\]\[1\] _01278_ _01942_ VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__mux2_1
X_09635_ _03350_ _03383_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06847_ _00964_ _00619_ _00629_ _00971_ VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__a211o_1
X_06778_ _00905_ VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__clkbuf_1
X_09566_ _03471_ _03474_ VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08517_ Oset\[2\]\[12\] VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__inv_2
X_09497_ _03380_ _03406_ VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08448_ _02356_ Oset\[1\]\[9\] _02329_ _02369_ VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__a211o_1
XFILLER_0_92_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10410_ _04313_ _04315_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__nand2_1
X_08379_ H\[1\]\[6\] _02260_ VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__nor2_1
X_11390_ _05289_ _05291_ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_21_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10341_ _04196_ _04246_ _04247_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__or3_2
XFILLER_0_33_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10272_ _03986_ _04160_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12011_ _05844_ _00658_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__nand2_1
X_12913_ clknet_leaf_15_clk _00356_ VGND VGND VPWR VPWR result_reg_or\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ clknet_leaf_8_clk _00287_ VGND VGND VPWR VPWR result_reg_mul\[11\] sky130_fd_sc_hd__dfxtp_1
X_12775_ clknet_leaf_27_clk _00218_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _05625_ VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11657_ _04189_ _04181_ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11588_ _05487_ _05488_ VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__nand2_1
X_10608_ _04512_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__inv_2
X_10539_ _02653_ _04444_ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12209_ _03846_ _04288_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__nand2_1
X_07750_ _01805_ _01589_ VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__nand2_1
X_06701_ _00536_ VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__clkbuf_4
X_07681_ _01740_ H\[3\]\[5\] _01629_ VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__mux2_1
X_06632_ result_reg_sub\[3\] _00541_ _00763_ VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__o21ai_1
X_09420_ _02273_ _02161_ VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06563_ CMD_load VGND VGND VPWR VPWR _00697_ sky130_fd_sc_hd__inv_2
X_09351_ _03254_ _03255_ _03261_ VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__nand3_1
XFILLER_0_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08302_ _02129_ VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__buf_6
X_09282_ _03192_ VGND VGND VPWR VPWR _03193_ sky130_fd_sc_hd__inv_2
X_06494_ _00628_ VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08233_ _02163_ _00591_ VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08164_ _02102_ _02103_ net39 VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__a21o_1
X_07115_ _01198_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__clkinv_4
X_08095_ _01761_ H\[1\]\[6\] _02057_ VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07046_ _01139_ VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08997_ _02906_ _02907_ _02908_ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__nand3_1
X_07948_ _01977_ VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__clkbuf_1
X_07879_ _01926_ _01663_ _01927_ _01928_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_54_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10890_ _04792_ _04793_ VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_26_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09618_ _03525_ _03526_ VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__nand2_1
X_09549_ _02821_ _03079_ VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12560_ _06214_ _05134_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__and2_1
X_12491_ _06211_ VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__clkbuf_1
X_11511_ _05225_ _05222_ VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__nand2_1
X_11442_ H\[2\]\[14\] _04856_ _05342_ VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11373_ _05104_ _05103_ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10324_ _04229_ _04230_ _03270_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__nand3_1
X_10255_ _04161_ _04149_ VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__nand2_1
X_10186_ _04090_ _04092_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_6_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12827_ clknet_leaf_12_clk _00270_ VGND VGND VPWR VPWR result_reg_sub\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12758_ clknet_leaf_53_clk _00201_ VGND VGND VPWR VPWR H\[0\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11709_ _01538_ _05608_ _00820_ VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12689_ clknet_leaf_52_clk _00139_ VGND VGND VPWR VPWR Oset\[0\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08920_ _02831_ _02832_ _00536_ VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__a21o_1
X_08851_ _02580_ Oset\[2\]\[2\] VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__nand2_1
X_07802_ _01716_ _01000_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__nand2_1
X_08782_ _02626_ _02693_ _02695_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__o21a_1
X_07733_ _01579_ result_reg_sub\[8\] VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07664_ _01722_ _01549_ _01723_ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__a21o_1
X_06615_ _00742_ _00743_ _00746_ _00747_ VGND VGND VPWR VPWR _00748_ sky130_fd_sc_hd__a31o_1
X_09403_ _03311_ _03312_ _03305_ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__nand3_1
XFILLER_0_94_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07595_ _01559_ VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06546_ R2\[0\] VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__inv_2
X_09334_ _02783_ _02213_ _02904_ VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__a21oi_1
X_06477_ _00610_ _00542_ _00611_ VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09265_ _03174_ _03175_ VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__nand2_2
XFILLER_0_7_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08216_ _02135_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_31_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09196_ _03080_ _03106_ VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__nand2_1
X_08147_ H\[0\]\[15\] _01938_ _02074_ VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08078_ _01938_ H\[2\]\[15\] _02037_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_591 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07029_ _00722_ Qset\[2\]\[1\] _01129_ VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__mux2_1
X_10040_ _03906_ _03946_ VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__xor2_1
X_11991_ result_reg_Lshift\[12\] _05741_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_3_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10942_ _03759_ Qset\[0\]\[12\] VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_11_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10873_ _04775_ _04593_ _04589_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__nand3b_1
X_12612_ clknet_leaf_43_clk _00062_ VGND VGND VPWR VPWR Qset\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_100_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12543_ _06242_ VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12474_ _06165_ _06129_ VGND VGND VPWR VPWR _06200_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_20_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11425_ _05319_ Qset\[3\]\[14\] _04303_ _05325_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__a211o_1
XANTENNA_7 _00621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11356_ _05095_ _05094_ _05099_ VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10307_ _04212_ _04201_ VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__nand2_1
X_13026_ clknet_leaf_54_clk _00469_ VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__dfxtp_2
X_11287_ _05187_ _05188_ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__nor2_1
X_10238_ _04111_ _04144_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__xor2_1
X_10169_ Qset\[1\]\[15\] VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06400_ _00534_ VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07380_ _00981_ _01275_ _01160_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06331_ _06285_ next_PC\[0\] VGND VGND VPWR VPWR _00476_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09050_ _02960_ _02961_ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08001_ Oset\[0\]\[11\] _01455_ _02000_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09952_ _03858_ VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__buf_6
XFILLER_0_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08903_ _02529_ _02207_ _02526_ _02815_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_57_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09883_ _03789_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__buf_6
X_08834_ _02744_ _02745_ _02747_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__a21o_1
X_08765_ _02579_ _02186_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__nor2_1
X_07716_ result_reg_mul\[7\] _01585_ _01589_ VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_0_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08696_ _02592_ VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__buf_6
X_07647_ _01581_ result_reg_add\[4\] VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07578_ _01586_ result_reg_sub\[1\] VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06529_ _00594_ _00661_ _00663_ VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__a21o_4
XFILLER_0_35_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09317_ _03218_ _03219_ _03227_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__nand3_2
XFILLER_0_90_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09248_ _03157_ Qset\[1\]\[4\] _02526_ _03158_ VGND VGND VPWR VPWR _03159_ sky130_fd_sc_hd__a211o_1
X_09179_ _02544_ Oset\[1\]\[6\] _02727_ _03089_ VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__a211o_1
XFILLER_0_16_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12190_ _03502_ _03102_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__nand2_1
X_11210_ _05055_ _05112_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_8_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11141_ _05029_ _05034_ _05033_ VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__a21bo_1
Xoutput44 net44 VGND VGND VPWR VPWR data_address[6] sky130_fd_sc_hd__buf_1
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput66 net66 VGND VGND VPWR VPWR instruction_address[1] sky130_fd_sc_hd__buf_1
Xoutput55 net55 VGND VGND VPWR VPWR data_out[1] sky130_fd_sc_hd__buf_1
XFILLER_0_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11072_ _04974_ _03079_ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__nand2_2
X_10023_ _02963_ _03876_ VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11974_ result_reg_Lshift\[9\] _05743_ _05808_ _05815_ VGND VGND VPWR VPWR _00317_
+ sky130_fd_sc_hd__o211a_1
X_10925_ _02654_ _04826_ _04828_ VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_62_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10856_ _04571_ _04568_ _04757_ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__nand3_1
XFILLER_0_39_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10787_ _04690_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_14_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12526_ _06232_ VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12457_ _06186_ _06117_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11408_ _05120_ _05129_ _05309_ VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_22_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12388_ _06123_ VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__inv_2
X_11339_ _05239_ _05240_ VGND VGND VPWR VPWR _05241_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06880_ _00998_ _01003_ VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__nand2_2
X_13009_ clknet_leaf_49_clk _00452_ VGND VGND VPWR VPWR Qset\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08550_ _02467_ _02444_ VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__nand2_1
X_07501_ _00569_ _01543_ VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__nand2_1
X_08481_ _02400_ _02397_ _02378_ _02401_ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07432_ _01499_ _01245_ _01502_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07363_ Oset\[3\]\[10\] _01437_ _01249_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__mux2_1
X_09102_ _02611_ H\[0\]\[4\] VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__nor2_1
X_07294_ net14 _01255_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__or2_1
X_06314_ LC\[3\] _06274_ VGND VGND VPWR VPWR _06275_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09033_ _02944_ _02572_ VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09935_ _03157_ _02368_ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__nor2_1
X_09866_ _03341_ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__buf_6
X_08817_ _02730_ _02571_ _00586_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__a21oi_1
X_09797_ _03682_ _03704_ _00624_ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__nand3_1
X_08748_ _02661_ _00580_ VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__nand2_1
X_08679_ _02589_ _02591_ _02593_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__nand3_1
XFILLER_0_95_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10710_ _04414_ H\[0\]\[10\] _03798_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11690_ _05556_ _05589_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10641_ _04042_ _04541_ _04543_ _04545_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_36_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10572_ _04474_ _04476_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__nand2_1
X_12311_ _06055_ _01390_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_11_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12242_ result_reg_or\[15\] _05960_ _06027_ _06029_ _02101_ VGND VGND VPWR VPWR _00371_
+ sky130_fd_sc_hd__o221a_1
X_12173_ _05969_ _05972_ _05957_ _04827_ _05973_ VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__o311a_1
X_11124_ _05010_ _05026_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11055_ _03790_ _04957_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__nand2_1
X_10006_ _03905_ _03912_ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_47_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ _05799_ _05766_ _05755_ _05800_ VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10908_ _01538_ _04811_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11888_ _05738_ _05739_ VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10839_ _04736_ _04742_ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12509_ next_PC\[2\] _06218_ VGND VGND VPWR VPWR _06224_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07981_ Oset\[0\]\[1\] _01278_ _02001_ VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__mux2_1
X_06932_ _01048_ _01053_ VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__nand2_2
X_09720_ _03498_ _02320_ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__nor2_1
X_06863_ result_reg_and\[11\] _00561_ _00553_ VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__o21ai_1
X_09651_ _03557_ _03559_ VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__nand2_1
X_06794_ _00654_ VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__inv_2
X_08602_ _02517_ _02444_ VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__nand2_1
X_09582_ _02295_ _02161_ VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08533_ _02451_ VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_85_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08464_ _02356_ _02384_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__nor2_1
X_07415_ _01486_ _01238_ _01215_ VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__o21ai_1
X_08395_ _02248_ VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__buf_4
XFILLER_0_18_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07346_ _01421_ VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07277_ _01353_ _01355_ _01181_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__mux2_1
X_09016_ _02586_ Qset\[3\]\[3\] VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09918_ _03824_ _02552_ VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__nand2_1
X_09849_ _03755_ _03752_ VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__nand2_1
X_12860_ clknet_leaf_10_clk _00303_ VGND VGND VPWR VPWR result_reg_mac\[11\] sky130_fd_sc_hd__dfxtp_2
X_11811_ _05686_ VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ clknet_leaf_45_clk _00234_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _00770_ _05631_ _05634_ _05637_ VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11673_ _05389_ _05380_ _05388_ VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_24_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10624_ _04157_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10555_ _03897_ _02897_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__nor2_1
X_10486_ _04364_ _04366_ _04391_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__nand3_1
XFILLER_0_32_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12225_ _04836_ _01666_ _05938_ VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__a21o_1
X_12156_ _05958_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11107_ _04919_ _04913_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__nand2_1
X_12087_ _03169_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_3_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11038_ _04923_ _04940_ VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12989_ clknet_leaf_7_clk _00432_ VGND VGND VPWR VPWR Oim sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07200_ result_reg_add\[2\] result_reg_sub\[2\] _01202_ VGND VGND VPWR VPWR _01283_
+ sky130_fd_sc_hd__mux2_1
X_08180_ _02095_ _02099_ net47 VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07131_ result_reg_mac\[0\] _01215_ VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07062_ _01148_ VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__buf_6
XFILLER_0_100_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07964_ im_reg\[7\] VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__inv_2
X_06915_ _01035_ _01036_ _00611_ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07895_ _01943_ VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__clkbuf_1
X_09703_ _03610_ VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__inv_2
X_06846_ _00965_ _00709_ _00603_ _00970_ VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__o211a_1
X_09634_ _03389_ _03384_ _03386_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__a21oi_1
X_06777_ _00904_ Qset\[0\]\[7\] _00687_ VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__mux2_1
X_09565_ _03473_ VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__inv_2
X_08516_ _02431_ _02434_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__nand2_2
X_09496_ _03404_ _03405_ VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__nand2_1
X_08447_ _02356_ _02368_ VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__nor2_1
X_08378_ H\[0\]\[6\] VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07329_ result_reg_Lshift\[9\] result_reg_Rshift\[9\] _01165_ VGND VGND VPWR VPWR
+ _01405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10340_ _04242_ _04244_ _04243_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__a21oi_1
X_10271_ _04172_ _04176_ _04177_ VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__a21oi_1
X_12010_ _02118_ _05759_ VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__nor2_1
X_12912_ clknet_leaf_16_clk _00355_ VGND VGND VPWR VPWR result_reg_and\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_57_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12843_ clknet_leaf_56_clk _00286_ VGND VGND VPWR VPWR result_reg_mul\[10\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12774_ clknet_leaf_28_clk _00217_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _05623_ _05624_ VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11656_ _05378_ _05398_ _05401_ VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__o21ai_1
X_11587_ result_reg_add\[14\] _02649_ _01149_ VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__o21a_1
X_10607_ _04510_ _04511_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10538_ _04442_ _04443_ VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__nand2_2
XFILLER_0_10_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12208_ _05960_ _06001_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__nand2_1
X_10469_ _04129_ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12139_ result_reg_and\[13\] _05894_ _05941_ _05944_ _05940_ VGND VGND VPWR VPWR
+ _00353_ sky130_fd_sc_hd__o221a_1
XFILLER_0_19_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06700_ _00528_ _00631_ _00634_ _00829_ VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__or4_1
X_07680_ _01736_ _01739_ _01613_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__mux2_4
X_06631_ _00740_ _00762_ _00535_ VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__a21oi_1
X_06562_ _00601_ VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__buf_2
XFILLER_0_87_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09350_ _03259_ VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__inv_2
X_08301_ _02225_ _02228_ VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__nand2_1
X_09281_ _03077_ _03190_ VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__nand2_1
X_06493_ _00620_ _00621_ _00625_ _00627_ VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__or4_4
X_08232_ _02162_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_62_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08163_ _01148_ VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__buf_4
XFILLER_0_27_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07114_ _01196_ _01198_ VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__nand2_4
X_08094_ _02063_ VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__clkbuf_1
X_07045_ _00953_ Qset\[2\]\[9\] _01129_ VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08996_ _02822_ _02899_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__nand2_1
X_07947_ _01976_ LC\[3\] _01964_ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07878_ result_reg_mul\[15\] _01688_ _01667_ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06829_ _00954_ VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_26_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09617_ _03519_ _03520_ _03523_ VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__nand3_1
X_09548_ _03453_ _03456_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11510_ _05409_ _05410_ _03746_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__nand3_2
X_09479_ _03387_ _03388_ VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12490_ _01151_ _05134_ VGND VGND VPWR VPWR _06211_ sky130_fd_sc_hd__and2_1
X_11441_ H\[3\]\[14\] _04858_ _04859_ VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11372_ _05272_ _05273_ VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10323_ _04226_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__inv_2
X_10254_ _04148_ _04146_ VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__or2_1
X_10185_ _03152_ H\[3\]\[15\] _02560_ _04091_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12826_ clknet_leaf_12_clk _00269_ VGND VGND VPWR VPWR result_reg_sub\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12757_ clknet_leaf_49_clk _00200_ VGND VGND VPWR VPWR H\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_11708_ _05603_ _05607_ _00647_ VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12688_ clknet_leaf_45_clk _00138_ VGND VGND VPWR VPWR Oset\[0\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11639_ _05537_ _03274_ _05536_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__nand3_1
XFILLER_0_12_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08850_ _02761_ _02762_ _02539_ VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__nand3_1
X_07801_ _01854_ result_reg_mac\[11\] _01540_ VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__mux2_1
X_08781_ Qset\[0\]\[1\] _02632_ _02694_ VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__a21o_1
X_07732_ _01580_ result_reg_add\[8\] VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__nand2_1
X_07663_ result_reg_mul\[5\] _01679_ _01561_ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06614_ result_reg_and\[2\] _00561_ _00552_ VGND VGND VPWR VPWR _00747_ sky130_fd_sc_hd__o21ai_2
X_09402_ _03245_ _03307_ VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__nand2_1
X_07594_ _00726_ _01656_ VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09333_ _03239_ _03242_ _03243_ VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__nand3_1
X_06545_ R0\[0\] _00602_ _00628_ VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__o21a_1
X_06476_ _00538_ _00574_ VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__nand2_4
X_09264_ _00498_ _00588_ VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09195_ _03104_ _03105_ VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__nand2_2
X_08215_ Oset\[0\]\[0\] VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08146_ _02090_ VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08077_ _02053_ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07028_ _01130_ VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__clkbuf_1
X_08979_ _02887_ _02888_ _02890_ VGND VGND VPWR VPWR _02891_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_97_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11990_ _05776_ _05817_ _02118_ _05828_ VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__o22a_1
X_10941_ _03759_ Qset\[2\]\[12\] _03345_ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_3_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12611_ clknet_leaf_45_clk _00061_ VGND VGND VPWR VPWR Qset\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_10872_ _04761_ _04775_ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_100_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12542_ _00904_ Qset\[3\]\[7\] _06234_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12473_ _06133_ _06149_ _06129_ _06139_ VGND VGND VPWR VPWR _06199_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11424_ _05319_ _02476_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__nor2_1
XANTENNA_8 _00626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11355_ _04281_ _05158_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__nor2_1
X_10306_ _04201_ _04212_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11286_ _04938_ _04935_ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__and2_1
X_13025_ clknet_leaf_52_clk _00468_ VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__dfxtp_2
X_10237_ _04114_ _04115_ _04113_ VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__o21ai_1
X_10168_ _04074_ _02620_ VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10099_ _04003_ _04005_ VGND VGND VPWR VPWR _04006_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12809_ clknet_leaf_10_clk _00252_ VGND VGND VPWR VPWR result_reg_add\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06330_ _00474_ VGND VGND VPWR VPWR _00475_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08000_ _02012_ VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09951_ _03856_ _03857_ VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__nand2_2
XFILLER_0_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08902_ _02545_ H\[3\]\[2\] VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__nand2_1
X_09882_ _03788_ _02353_ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__nand2_2
X_08833_ _02746_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__inv_2
X_08764_ _02585_ H\[1\]\[1\] _00005_ _02677_ VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__a211o_1
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07715_ _01586_ result_reg_sub\[7\] VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_88_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08695_ _02608_ _02609_ VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__nand2_1
X_07646_ _01704_ _01635_ _01705_ _01706_ VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07577_ _01581_ result_reg_add\[1\] VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__nand2_1
X_06528_ _00595_ CMD_not _00662_ VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__and3_1
X_09316_ _03226_ VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09247_ _02544_ Qset\[0\]\[4\] VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__and2b_1
XFILLER_0_90_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06459_ _00593_ _00531_ VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09178_ _02874_ _02299_ VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08129_ H\[0\]\[6\] _01761_ _02075_ VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__mux2_1
X_11140_ _05042_ _05038_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_8_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput45 net45 VGND VGND VPWR VPWR data_address[7] sky130_fd_sc_hd__buf_1
Xoutput56 net56 VGND VGND VPWR VPWR data_out[2] sky130_fd_sc_hd__buf_1
Xoutput67 net67 VGND VGND VPWR VPWR instruction_address[2] sky130_fd_sc_hd__buf_1
X_11071_ _04973_ VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__inv_2
X_10022_ _03879_ _03928_ VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11973_ _05814_ _05771_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__nand2_1
X_10924_ result_reg_add\[11\] _02649_ _04827_ VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_62_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10855_ _04724_ _04758_ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12525_ _00685_ _01126_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_70_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10786_ _04689_ _02426_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__nand2_8
XTAP_TAPCELL_ROW_42_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12456_ _06132_ _06128_ VGND VGND VPWR VPWR _06186_ sky130_fd_sc_hd__nand2_1
X_12387_ _06128_ _06256_ VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__nand2_1
X_11407_ _05117_ _03296_ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__and2_1
X_11338_ _05238_ _05234_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11269_ _04855_ H\[0\]\[13\] _04862_ VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__a21oi_1
X_13008_ clknet_leaf_34_clk _00451_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dfxtp_1
X_07500_ _01550_ _01562_ _01563_ _01564_ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__a211o_1
X_08480_ _02397_ H\[0\]\[10\] VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__nor2_1
X_07431_ _01060_ _01265_ _01206_ _01501_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07362_ _01276_ _01423_ _01435_ _01436_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__a22o_2
XFILLER_0_91_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06313_ LC\[2\] _06273_ VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09101_ _02611_ H\[2\]\[4\] _02584_ VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__o21ai_1
X_07293_ result_reg_not\[7\] _01370_ _01168_ VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09032_ _02943_ VGND VGND VPWR VPWR _02944_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09934_ _02162_ _03840_ _02713_ VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09865_ _03759_ Oset\[0\]\[8\] VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__nor2_1
X_08816_ _02726_ _02727_ _02728_ _02729_ VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__a22oi_4
X_09796_ _03701_ _03703_ _03233_ VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__nand3_2
X_08747_ _02657_ _02660_ VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__nand2_2
X_08678_ Qset\[1\]\[0\] _02592_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__nand2_1
X_07629_ _01577_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10640_ _04105_ Oset\[3\]\[10\] _04045_ _04544_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10571_ _04282_ Qset\[1\]\[10\] _03345_ _04475_ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__a211o_1
XFILLER_0_36_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12310_ _05766_ _01959_ _03834_ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_11_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12241_ _05904_ _05515_ _06028_ _00524_ _05951_ VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12172_ _05957_ _00738_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11123_ _05024_ _05025_ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__and2_1
X_11054_ _04956_ VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__inv_2
X_10005_ _03907_ _03910_ _03911_ VGND VGND VPWR VPWR _03912_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_47_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ _05755_ _05785_ VGND VGND VPWR VPWR _05800_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10907_ _04805_ _04810_ _00621_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__mux2_1
X_11887_ result_reg_mac\[15\] _05703_ _01149_ VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10838_ _02163_ _04741_ _02872_ VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10769_ _04282_ _02406_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12508_ net66 _06220_ _06221_ _06223_ VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__o211a_1
X_12439_ _06171_ _06157_ _06172_ _06106_ VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07980_ _02002_ VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__clkbuf_1
X_06931_ _01049_ _00654_ _00656_ _01052_ _00665_ VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__a221o_1
X_09650_ _03558_ _03556_ _03554_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__nand3_1
X_06862_ _00985_ _00745_ VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__or2_1
X_08601_ H\[2\]\[15\] H\[3\]\[15\] _02491_ VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__mux2_1
X_06793_ _00695_ _00919_ VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__nand2_1
X_09581_ _03489_ _00581_ VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__nand2_1
X_08532_ _02450_ net51 _02169_ VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08463_ Oset\[2\]\[10\] VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__inv_2
X_07414_ _01482_ _01485_ _01041_ _01271_ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_64_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08394_ _02314_ _02317_ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__nand2_2
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07345_ Oset\[3\]\[9\] _01420_ _01250_ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__mux2_1
X_07276_ _00860_ _01354_ _01176_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_30_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09015_ _02582_ Qset\[2\]\[3\] VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_96_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09917_ _03821_ _03822_ _03823_ _02560_ VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__a22oi_4
X_09848_ _03750_ _03746_ _03744_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__nand3_1
X_09779_ _03507_ _03383_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__nor2_1
X_11810_ _03682_ _03704_ _05677_ _05685_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__a31o_1
X_12790_ clknet_leaf_45_clk _00233_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dfxtp_1
X_11741_ _05631_ _02986_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11672_ _05570_ _05571_ VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_24_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10623_ _04398_ _04192_ _04159_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_21_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
X_10554_ _04458_ _04309_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10485_ _04387_ _04390_ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__nand2_1
X_12224_ _04891_ _04847_ _05892_ VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__a21oi_1
X_12155_ _05957_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__inv_2
X_11106_ _05007_ _05008_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__and2_1
X_12086_ _05767_ _00524_ _02994_ _02997_ _05872_ VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__a41o_1
X_11037_ _04938_ _04939_ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12988_ clknet_leaf_0_clk _00431_ VGND VGND VPWR VPWR Oreg3 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_24_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11939_ _05744_ _05783_ _05784_ VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__a21o_2
XFILLER_0_74_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07130_ _01214_ VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_12_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07061_ _00472_ VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07963_ _01986_ _01987_ _01989_ LC\[6\] VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__a22o_1
X_06914_ result_reg_add\[13\] VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__inv_2
X_07894_ Oset\[2\]\[0\] _01218_ _01942_ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__mux2_1
X_09702_ _03465_ _03461_ _03609_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__a21oi_2
X_06845_ _00967_ _00743_ _00968_ _00969_ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09633_ _03507_ _03206_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__nor2_1
X_09564_ _03306_ _03309_ _03472_ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__a21oi_2
X_06776_ _00664_ _00898_ _00903_ VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__o21ai_4
X_08515_ _02328_ Qset\[1\]\[12\] _02329_ _02433_ VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__a211o_1
XFILLER_0_77_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09495_ _03381_ _03402_ _03401_ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__nand3_1
X_08446_ Oset\[0\]\[9\] VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08377_ _02298_ _02301_ VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_98_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07328_ _01404_ VGND VGND VPWR VPWR _00082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07259_ net12 _01193_ VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10270_ _04171_ _04169_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__nor2_1
X_12911_ clknet_leaf_17_clk _00354_ VGND VGND VPWR VPWR result_reg_and\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_57_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ clknet_leaf_56_clk _00285_ VGND VGND VPWR VPWR result_reg_mul\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_96_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12773_ clknet_leaf_27_clk _00216_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ result_reg_add\[15\] _02649_ _01149_ VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__o21a_1
X_11655_ _05409_ _05405_ VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11586_ _05485_ _02649_ _05486_ VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__nand3_1
XFILLER_0_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10606_ _03564_ _04507_ _04508_ VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__nand3b_1
X_10537_ _04441_ _04255_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10468_ _04125_ _04097_ VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__nor2_1
X_12207_ _04294_ _03840_ _05907_ VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_71_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10399_ _03764_ _04300_ _04301_ _04304_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__o2bb2a_1
X_12138_ _05825_ _05942_ _05943_ _05154_ VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__a22o_1
X_12069_ _05883_ _05885_ _05886_ _05878_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_1_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
X_06630_ result_reg_add\[3\] VGND VGND VPWR VPWR _00762_ sky130_fd_sc_hd__inv_2
X_06561_ _00650_ VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_82_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06492_ _00472_ _00626_ VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__nand2_1
X_08300_ _02141_ _02226_ _02147_ _02227_ VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__o211ai_1
X_09280_ _03077_ _03190_ VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08231_ _02161_ VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__clkbuf_4
X_08162_ R3\[0\] _02100_ _02101_ _02104_ VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07113_ Hreg2 _01197_ VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__nor2_4
X_08093_ _01740_ H\[1\]\[5\] _02057_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__mux2_1
X_07044_ _01138_ VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_93_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08995_ _02901_ VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07946_ _01960_ _00671_ _01975_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__a21oi_1
X_07877_ _01579_ result_reg_sub\[15\] VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__nand2_1
X_06828_ _00953_ Qset\[0\]\[9\] _00687_ VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__mux2_1
X_09616_ _03521_ _03524_ VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__nand2_1
X_06759_ _00881_ _00886_ _00608_ VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09547_ _03264_ _03454_ _03455_ VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__a21oi_1
X_09478_ _03116_ _03076_ VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_419 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08429_ _02327_ _02350_ _02329_ _02351_ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11440_ _05340_ _02497_ VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__nand2_4
XFILLER_0_33_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11371_ _05270_ _05256_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10322_ _03364_ _03266_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10253_ _03957_ _03984_ _03960_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__nand3_1
X_10184_ _02529_ H\[2\]\[15\] VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_6_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12825_ clknet_leaf_10_clk _00268_ VGND VGND VPWR VPWR result_reg_sub\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12756_ clknet_leaf_30_clk _00199_ VGND VGND VPWR VPWR H\[1\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11707_ _05604_ _05605_ _05606_ _04859_ VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__a22o_1
X_12687_ clknet_leaf_53_clk _00137_ VGND VGND VPWR VPWR Oset\[0\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11638_ _05536_ _05537_ _03274_ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11569_ _05411_ _05469_ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07800_ _01594_ _01846_ _01853_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__o21ai_1
X_08780_ Qset\[1\]\[1\] _02624_ _00001_ VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__a21o_1
X_07731_ _01785_ _01635_ _01786_ _01787_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__a31o_1
X_07662_ _00841_ _00812_ _01545_ VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06613_ _00727_ _00745_ VGND VGND VPWR VPWR _00746_ sky130_fd_sc_hd__or2_1
X_07593_ _01560_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__buf_2
X_09401_ _03308_ _02821_ _02963_ VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__nand3_1
X_06544_ _00678_ VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09332_ _02963_ _02734_ VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__nand2_1
X_06475_ result_reg_sub\[0\] VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__inv_2
X_09263_ _03156_ _03173_ VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09194_ _00587_ im_reg\[6\] VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__nand2_1
X_08214_ _02141_ _02142_ _02143_ _02144_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08145_ H\[0\]\[14\] _01918_ _02074_ VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08076_ _01918_ H\[2\]\[14\] _02037_ VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__mux2_1
X_07027_ _00668_ Qset\[2\]\[0\] _01129_ VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08978_ _02798_ _02231_ _02525_ _02889_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_98_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07929_ CMD_setloop VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10940_ Qset\[3\]\[12\] _03773_ VGND VGND VPWR VPWR _04843_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_3_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10871_ _04762_ _04774_ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__xor2_1
X_12610_ clknet_leaf_48_clk _00060_ VGND VGND VPWR VPWR Qset\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12541_ _06241_ VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__clkbuf_1
X_12472_ _06097_ Oim _04827_ _06194_ VGND VGND VPWR VPWR _00432_ sky130_fd_sc_hd__o211a_1
X_11423_ _05321_ _05323_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_9 _00648_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11354_ _05101_ _05090_ _05255_ VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10305_ _04210_ _04211_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11285_ _05176_ _05186_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__xnor2_1
X_13024_ clknet_leaf_25_clk _00467_ VGND VGND VPWR VPWR Qset\[3\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_10236_ _04117_ _04119_ _04118_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__nand3_1
X_10167_ _02556_ _04073_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__nor2_4
XFILLER_0_83_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10098_ _04004_ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12808_ clknet_leaf_12_clk _00251_ VGND VGND VPWR VPWR result_reg_add\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12739_ clknet_leaf_25_clk _00182_ VGND VGND VPWR VPWR H\[2\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09950_ _00588_ im_reg\[9\] VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08901_ _02798_ H\[1\]\[2\] _02525_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09881_ _03787_ _01553_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__nand2_1
X_08832_ _00536_ _02643_ _02622_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__mux2_1
X_08763_ _02579_ _02189_ VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__nor2_1
X_07714_ _01581_ result_reg_add\[7\] VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08694_ _02150_ _00583_ _02571_ VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_36_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07645_ net11 _01658_ VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07576_ net8 _01635_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06527_ _00545_ VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__inv_2
X_09315_ _03223_ _03225_ VGND VGND VPWR VPWR _03226_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06458_ _00592_ VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09246_ _02798_ VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__buf_4
XFILLER_0_35_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06389_ Oreg2 Hreg2 VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__nor2_4
XFILLER_0_7_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09177_ _02544_ Oset\[3\]\[6\] _02534_ _03087_ VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__a211o_1
X_08128_ _02081_ VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08059_ _02044_ VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__clkbuf_1
Xoutput46 net46 VGND VGND VPWR VPWR data_address[8] sky130_fd_sc_hd__buf_1
X_11070_ _04971_ _04972_ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__nand2_1
Xoutput57 net57 VGND VGND VPWR VPWR data_out[3] sky130_fd_sc_hd__buf_1
Xoutput68 net68 VGND VGND VPWR VPWR instruction_address[3] sky130_fd_sc_hd__buf_1
X_10021_ _02963_ _03868_ VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11972_ _05812_ _05813_ _02118_ VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10923_ _00472_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10854_ _04757_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_70_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12524_ net74 _06220_ _06221_ _06231_ VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__o211a_1
X_10785_ _04688_ _01553_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_42_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12455_ _06139_ _06181_ _06123_ _06175_ VGND VGND VPWR VPWR _06185_ sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_3_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_12386_ net22 _06100_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__nor2_2
X_11406_ _05307_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11337_ _05234_ _05238_ VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11268_ H\[2\]\[13\] _04855_ _05169_ VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__a21o_1
X_13007_ clknet_leaf_35_clk _00450_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dfxtp_1
X_11199_ _05090_ _05101_ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__xnor2_1
X_10219_ _04097_ _04125_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07430_ _01067_ _01202_ _01204_ _01500_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07361_ _00955_ _01275_ _01160_ VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06312_ LC\[1\] LC\[0\] VGND VGND VPWR VPWR _06273_ sky130_fd_sc_hd__or2_1
X_09100_ H\[3\]\[4\] _02582_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__nor2_1
X_07292_ result_reg_Lshift\[7\] result_reg_Rshift\[7\] _01165_ VGND VGND VPWR VPWR
+ _01370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09031_ _02940_ _02942_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09933_ _03836_ _03837_ _03838_ _03839_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__o22a_4
XFILLER_0_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09864_ Oset\[2\]\[8\] Oset\[3\]\[8\] _03498_ VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__mux2_1
X_08815_ _02522_ _02189_ VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09795_ _03562_ _03702_ _03559_ VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__nand3_1
X_08746_ _02658_ _02590_ _02659_ VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__nand3_1
X_08677_ _02579_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__buf_6
X_07628_ _01686_ _01663_ _01687_ _01689_ VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07559_ _00681_ _01568_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10570_ _03759_ _02391_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__nor2_1
X_09229_ _03136_ H\[2\]\[5\] _03139_ VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__a21oi_1
X_12240_ _05836_ _05506_ VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__or2_1
X_12171_ _01243_ _05970_ _05971_ _01666_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11122_ _05022_ _05021_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__nand2_1
X_11053_ _04955_ _03079_ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10004_ _03887_ _03909_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11955_ _05796_ _05797_ _05798_ VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_47_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10906_ _04806_ _04807_ _03795_ _04808_ _04809_ VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__a32o_1
X_11886_ _05621_ _05622_ _05703_ VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_17_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10837_ _04738_ _04740_ VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__nand2_2
XFILLER_0_66_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10768_ _02412_ _02162_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__nand2_1
X_12507_ next_PC\[1\] _06218_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__or2_1
X_12438_ _06164_ _06128_ VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10699_ _04573_ _03751_ _03745_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12369_ net22 VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_26_Left_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06930_ result_reg_Rshift\[13\] _00753_ _01051_ VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06861_ result_reg_mul\[11\] VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__inv_2
X_08600_ _02327_ _02514_ _02444_ _02515_ VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__a211o_1
X_06792_ result_reg_mac\[8\] VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__inv_2
X_09580_ _03485_ _03486_ _03488_ VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__o21ai_2
X_08531_ _02311_ _02435_ _02139_ _02442_ _02449_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__o221ai_4
XTAP_TAPCELL_ROW_85_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08462_ _02383_ VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_35_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07413_ result_reg_mul\[13\] _01263_ _01245_ _01484_ VGND VGND VPWR VPWR _01485_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08393_ _02248_ Qset\[1\]\[7\] _02143_ _02316_ VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__a211o_1
X_07344_ _01161_ _01406_ _01419_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__a21bo_4
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07275_ _00865_ _00857_ _01173_ VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09014_ _02222_ _02161_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_44_Left_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09916_ Oset\[2\]\[8\] Oset\[3\]\[8\] _02798_ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__mux2_1
X_09847_ _03748_ _03750_ _03753_ VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__nand3_1
X_09778_ _03206_ _03685_ VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08729_ _00832_ _02643_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__xor2_2
X_11740_ _05636_ VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _05377_ _05375_ _05374_ VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_36_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10622_ _04525_ _03746_ _04526_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__nand3_2
XFILLER_0_8_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10553_ _04270_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_24_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10484_ _04388_ _04389_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__nand2_1
X_12223_ _04886_ _04842_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__or2_1
X_12154_ _05956_ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__clkbuf_4
X_11105_ _05006_ _04993_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__nand2_1
X_12085_ result_reg_and\[3\] _05894_ _05896_ _05900_ _02125_ VGND VGND VPWR VPWR _00343_
+ sky130_fd_sc_hd__o221a_1
X_11036_ _04924_ _04926_ _04937_ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12987_ clknet_leaf_6_clk _00430_ VGND VGND VPWR VPWR Oreg2 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11938_ _01158_ _03091_ _03102_ _05749_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__a22o_1
X_11869_ _05726_ VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07060_ R0\[0\] net18 _01146_ VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07962_ _01986_ _01988_ VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__nand2_1
X_09701_ _03464_ _03463_ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__nor2_1
X_06913_ result_reg_sub\[13\] VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__inv_2
X_07893_ _01941_ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__buf_4
X_06844_ result_reg_and\[10\] _00561_ _00552_ VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__o21ai_1
X_09632_ _03537_ _03540_ VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__nand2_1
X_09563_ _03238_ _03464_ VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__nor2_1
X_06775_ _00899_ _00655_ _00657_ _00902_ _00666_ VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__a221o_1
X_08514_ _02319_ _02432_ VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__nor2_1
X_09494_ _03382_ _03403_ VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08445_ _02364_ Oset\[3\]\[9\] _02347_ _02366_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__a211o_1
X_08376_ _02261_ Oset\[1\]\[6\] _02250_ _02300_ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__a211o_1
XFILLER_0_18_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07327_ Oset\[3\]\[8\] _01403_ _01250_ VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07258_ _00840_ _01337_ _01181_ VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07189_ _01272_ _01238_ _01215_ VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12910_ clknet_leaf_16_clk _00353_ VGND VGND VPWR VPWR result_reg_and\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_57_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12841_ clknet_leaf_56_clk _00284_ VGND VGND VPWR VPWR result_reg_mul\[8\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_29_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12772_ clknet_leaf_26_clk _00215_ VGND VGND VPWR VPWR H\[0\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _05621_ _02649_ _05622_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__nand3_1
X_11654_ _05531_ _05553_ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__nand2_1
X_10605_ _04509_ _03564_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11585_ _05484_ _05483_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10536_ _04255_ _04441_ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10467_ _04371_ _04372_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__nand2_1
X_12206_ result_reg_or\[8\] _05959_ _05997_ _06000_ _05940_ VGND VGND VPWR VPWR _00364_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10398_ H\[1\]\[9\] _04302_ _04303_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__o21ai_1
X_12137_ _05888_ _04047_ VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__nor2_1
X_12068_ _00525_ _02711_ _02661_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__or3_1
X_11019_ _04568_ _04757_ _04755_ VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06560_ result_reg_mac\[1\] VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06491_ Hreg3 VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__inv_4
XFILLER_0_47_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08230_ shift.Q VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08161_ _02102_ _02103_ net38 VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07112_ Oreg2 VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__inv_2
X_08092_ _02062_ VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07043_ _00927_ Qset\[2\]\[8\] _01129_ VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08994_ _02903_ _02905_ VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__nand2_1
X_07945_ _06275_ _01962_ _01974_ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__and3_1
X_07876_ _01580_ result_reg_add\[15\] VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__nand2_1
X_09615_ _03523_ VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__inv_2
X_06827_ _00664_ _00947_ _00952_ VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__o21ai_4
X_06758_ _00882_ _00885_ _00732_ VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09546_ _03357_ _03354_ VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09477_ _03184_ _03110_ VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__nand2_1
X_06689_ _00714_ result_reg_or\[5\] VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08428_ H\[1\]\[8\] _02327_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08359_ _02260_ H\[3\]\[5\] _02284_ VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__o21ai_1
X_11370_ _05271_ VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10321_ _04225_ _04227_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10252_ _04158_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__inv_2
X_10183_ H\[1\]\[15\] _03152_ _03135_ _04089_ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_6_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12824_ clknet_leaf_12_clk _00267_ VGND VGND VPWR VPWR result_reg_sub\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12755_ clknet_leaf_26_clk _00198_ VGND VGND VPWR VPWR H\[1\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_11706_ _02503_ _04076_ _03793_ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12686_ clknet_leaf_53_clk _00136_ VGND VGND VPWR VPWR Oset\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11637_ _04607_ _05158_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__nor2_1
X_11568_ _05468_ _04196_ VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10519_ Oset\[3\]\[9\] _03791_ _03794_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11499_ _05359_ _05399_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_20_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07730_ net15 _01746_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07661_ _01721_ VGND VGND VPWR VPWR _00098_ sky130_fd_sc_hd__clkbuf_1
X_07592_ _01652_ _01549_ _01654_ VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06612_ _00744_ VGND VGND VPWR VPWR _00745_ sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_9_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09400_ _03302_ _03306_ _03309_ VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__nand3_1
X_06543_ _00675_ _00677_ VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__nand2_1
X_09331_ _03240_ _03241_ VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06474_ result_reg_mul\[0\] VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__inv_2
X_09262_ _03171_ _02556_ _03172_ VGND VGND VPWR VPWR _03173_ sky130_fd_sc_hd__nand3_1
XFILLER_0_90_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09193_ _03097_ _03103_ VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__nand2_1
X_08213_ _02141_ Oset\[3\]\[0\] VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08144_ _02089_ VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_31_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08075_ _02052_ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07026_ _01128_ VGND VGND VPWR VPWR _01129_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_87_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08977_ _02798_ H\[3\]\[3\] VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__nand2_1
X_07928_ LC\[0\] _01959_ _01960_ VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07859_ _01691_ result_reg_and\[14\] VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10870_ _04763_ _04773_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09529_ _00623_ _03421_ _03438_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_100_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12540_ _00878_ Qset\[3\]\[6\] _06234_ VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12471_ _02116_ _06198_ VGND VGND VPWR VPWR _00431_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11422_ _05319_ Oset\[1\]\[14\] _04835_ _05322_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11353_ _05091_ _05100_ VGND VGND VPWR VPWR _05255_ sky130_fd_sc_hd__nor2_1
X_10304_ _04203_ _04206_ _04208_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11284_ _05184_ _05185_ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__and2b_1
X_13023_ clknet_leaf_25_clk _00466_ VGND VGND VPWR VPWR Qset\[3\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_10235_ _02949_ _04110_ _04141_ VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__o21ai_1
X_10166_ _04066_ _04072_ VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__nand2_4
X_10097_ _03978_ _03972_ VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12807_ clknet_leaf_11_clk _00250_ VGND VGND VPWR VPWR result_reg_add\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10999_ _04074_ _03506_ _04096_ _03421_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__a22o_1
X_12738_ clknet_leaf_25_clk _00181_ VGND VGND VPWR VPWR H\[2\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12669_ clknet_leaf_40_clk _00119_ VGND VGND VPWR VPWR Oset\[2\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08900_ _02529_ _02210_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__nor2_1
X_09880_ _03758_ _03767_ _03769_ _03786_ VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__o22ai_1
X_08831_ _02743_ _02704_ VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__nand2_1
X_08762_ _02674_ _02675_ VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__nand2_1
X_07713_ _01768_ _01635_ _01769_ _01593_ _01770_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__a311o_1
X_08693_ _02598_ _02607_ VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__nand2_1
X_07644_ _00786_ _01682_ VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07575_ _00700_ _01561_ _01635_ _01638_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_48_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06526_ _00546_ _00639_ VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__nor2_2
X_09314_ _03179_ _03224_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__nor2_1
X_06457_ _00582_ _00591_ VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__nor2_2
X_09245_ _03155_ _02573_ _00588_ VGND VGND VPWR VPWR _03156_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06388_ Qreg2 VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__inv_2
X_09176_ _02874_ _02296_ VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08127_ H\[0\]\[5\] _01740_ _02075_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08058_ _01740_ H\[2\]\[5\] _02038_ VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__mux2_1
Xoutput47 net47 VGND VGND VPWR VPWR data_address[9] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_8_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07009_ _00953_ Qset\[1\]\[9\] _01109_ VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__mux2_1
Xoutput36 net36 VGND VGND VPWR VPWR data_R sky130_fd_sc_hd__buf_1
Xoutput58 net58 VGND VGND VPWR VPWR data_out[4] sky130_fd_sc_hd__buf_1
XFILLER_0_31_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput69 net69 VGND VGND VPWR VPWR instruction_address[4] sky130_fd_sc_hd__buf_1
X_10020_ _03858_ _03050_ _03020_ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__nand3_1
X_11971_ _05799_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__inv_2
X_10922_ _04824_ _04825_ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__xor2_2
XFILLER_0_85_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10853_ _04755_ _04756_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__nand2_2
XFILLER_0_66_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10784_ _03768_ _04671_ _04686_ _04687_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__a22o_1
X_12523_ next_PC\[9\] _06218_ VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12454_ _06177_ _06184_ _02650_ VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__a21oi_1
X_12385_ _06125_ _06127_ _02116_ VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__a21oi_1
X_11405_ _05303_ _05306_ VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__nand2_1
X_11336_ _05067_ _05235_ _05237_ VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__o21a_1
X_11267_ H\[3\]\[13\] _04857_ _04859_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__a21o_1
X_13006_ clknet_leaf_35_clk _00449_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dfxtp_1
X_11198_ _05091_ _05100_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__xor2_1
X_10218_ _04074_ _02785_ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__nand2_1
X_10149_ _03157_ Qset\[3\]\[14\] _02535_ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_99_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07360_ _01254_ _01424_ _01428_ _01434_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06311_ _06272_ VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07291_ _01369_ VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09030_ _02592_ H\[1\]\[3\] _00005_ _02941_ VGND VGND VPWR VPWR _02942_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09932_ Qset\[1\]\[9\] _03136_ _03135_ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__o21ai_1
X_09863_ _02540_ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__buf_4
X_08814_ H\[1\]\[1\] _02522_ _02534_ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__o21a_1
X_09794_ _03699_ _03700_ VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08745_ _02585_ Qset\[1\]\[1\] VGND VGND VPWR VPWR _02659_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08676_ _02590_ VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__buf_4
X_07627_ result_reg_mul\[3\] _01688_ _01667_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07558_ _01619_ _01622_ VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__or2b_1
X_06509_ _00633_ _00636_ _00594_ _00640_ _00643_ VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__a221o_4
XFILLER_0_63_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07489_ _01553_ VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__buf_4
X_09228_ _02798_ H\[3\]\[5\] _02800_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09159_ H\[1\]\[7\] _02522_ _02800_ VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__o21a_1
X_12170_ _02781_ _02817_ VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__nand2_1
X_11121_ _05023_ VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11052_ _04073_ VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__inv_2
X_10003_ _03909_ _03887_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11954_ _03831_ _00589_ VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_47_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11885_ _05737_ VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10905_ _04414_ Oset\[2\]\[11\] VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10836_ _04729_ Qset\[1\]\[11\] _04042_ _04739_ VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__a211o_1
XFILLER_0_13_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10767_ _04668_ _04669_ _04670_ _03764_ VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12506_ net65 _06220_ _06221_ _06222_ VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__o211a_1
X_10698_ _04602_ _03048_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12437_ _06170_ VGND VGND VPWR VPWR _06171_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12368_ _06112_ VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_74_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12299_ result_reg_set\[4\] _06063_ _06044_ _06065_ VGND VGND VPWR VPWR _00392_ sky130_fd_sc_hd__o211a_1
X_11319_ _05001_ _05004_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06860_ result_reg_sub\[11\] _00541_ _00983_ VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__o21ai_1
X_06791_ _00909_ _00910_ _00917_ _00619_ _00629_ VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__a221o_1
X_08530_ _02445_ _02448_ _01553_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_85_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08461_ _02382_ net63 _02170_ VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__mux2_1
X_07412_ result_reg_add\[13\] _01264_ _01266_ _01483_ VGND VGND VPWR VPWR _01484_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08392_ _02241_ _02315_ VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__nor2_1
X_07343_ _00929_ _01220_ _01160_ _01418_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__a211o_1
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07274_ result_reg_set\[6\] VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09013_ _02924_ VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09915_ Oset\[1\]\[8\] _02523_ _02535_ VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__o21a_1
X_09846_ _03752_ VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__inv_2
X_06989_ _00679_ _00684_ VGND VGND VPWR VPWR _01108_ sky130_fd_sc_hd__nand2_4
X_09777_ _03651_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__inv_2
X_08728_ _00622_ _02620_ _02642_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_68_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _02570_ _02573_ _00587_ VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_105_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11670_ _05559_ _05569_ VGND VGND VPWR VPWR _05570_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_52_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10621_ _04447_ _04523_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_24_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10552_ _04311_ _04456_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12222_ _01148_ VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10483_ _04153_ _04139_ _04138_ VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12153_ _00662_ _00572_ _05955_ _02167_ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__or4_1
X_12084_ _05897_ _05899_ VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__nand2_1
X_11104_ _04993_ _05006_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__or2_1
X_11035_ _04924_ _04926_ _04937_ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__or3_1
XFILLER_0_99_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12986_ clknet_leaf_5_clk _00429_ VGND VGND VPWR VPWR shift.O sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11937_ _03082_ _03084_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__nand2_1
X_11868_ _00929_ _05707_ _05710_ _05725_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__a211o_1
X_11799_ result_reg_mul\[4\] _05677_ _05134_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10819_ _04600_ _04597_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07961_ _01962_ im_reg\[6\] _06279_ VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__o21ai_1
X_06912_ result_reg_mul\[13\] VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09700_ _03519_ _03607_ VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__nand2_1
X_07892_ _01940_ _01248_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__nor2_4
X_06843_ _00957_ _00744_ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__or2_1
X_09631_ _03538_ _03214_ _03539_ VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__a21oi_1
X_06774_ _00900_ _00901_ _00643_ VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__mux2_1
X_09562_ _03466_ _03470_ VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08513_ Qset\[0\]\[12\] VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__inv_2
X_09493_ _03401_ _03402_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08444_ _02356_ _02365_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__nor2_1
X_08375_ _02248_ _02299_ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_98_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07326_ _01276_ _01388_ _01401_ _01402_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__a22o_4
XFILLER_0_73_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07257_ _00815_ _01336_ _01176_ VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07188_ _01262_ _01270_ _00708_ _01271_ VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__o2bb2a_1
X_09829_ _03735_ _03736_ VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_57_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12840_ clknet_leaf_56_clk _00283_ VGND VGND VPWR VPWR result_reg_mul\[7\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_29_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ clknet_leaf_26_clk _00214_ VGND VGND VPWR VPWR H\[0\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11722_ _05491_ _05482_ _05619_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__nand3_1
XFILLER_0_68_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11653_ _03751_ _05552_ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__or2_1
X_10604_ _04507_ _04508_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11584_ _05483_ _05484_ VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__or2_1
X_10535_ _04438_ _04440_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10466_ _04370_ _04368_ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12205_ _05904_ _05998_ _05999_ _05937_ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12136_ _05881_ _05141_ VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__nor2_1
X_10397_ _03761_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_63_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12067_ _05884_ _02682_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__nand2_1
X_11018_ _04757_ _04571_ VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__or2_1
X_12969_ clknet_leaf_7_clk _00412_ VGND VGND VPWR VPWR CMD_multiplication sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06490_ _00558_ _00624_ VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__nand2_2
XFILLER_0_59_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_72_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08160_ _02099_ VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__buf_2
XFILLER_0_51_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07111_ _00550_ _00471_ _00545_ _00558_ VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__and4_2
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08091_ _01720_ H\[1\]\[4\] _02057_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07042_ _01137_ VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_81_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08993_ _02685_ _02192_ _02904_ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__a21oi_1
X_07944_ _06274_ LC\[3\] VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__nand2_1
X_07875_ _01922_ _01658_ _01923_ _01924_ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06826_ _00948_ _00655_ _00657_ _00951_ _00666_ VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__a221o_1
X_09614_ _03522_ _03226_ VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__nand2_1
X_06757_ _00883_ _00884_ _00730_ VGND VGND VPWR VPWR _00885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09545_ _03354_ _03357_ VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__nand2_1
X_06688_ _00814_ _00562_ _00816_ _00817_ VGND VGND VPWR VPWR _00818_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_90_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09476_ _03190_ _03385_ VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__nor2_1
X_08427_ H\[0\]\[8\] VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_579 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08358_ _02261_ H\[2\]\[5\] _02250_ VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07309_ _01386_ VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08289_ _02131_ Qset\[3\]\[3\] VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__nand2_1
X_10320_ _04226_ _03456_ VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10251_ _04156_ _04157_ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__nand2_1
X_10182_ _03152_ _02514_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_6_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12823_ clknet_leaf_11_clk _00266_ VGND VGND VPWR VPWR result_reg_sub\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12754_ clknet_leaf_26_clk _00197_ VGND VGND VPWR VPWR H\[1\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_587 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11705_ Qset\[3\]\[15\] _04857_ _03795_ VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12685_ clknet_leaf_1_clk _00135_ VGND VGND VPWR VPWR LC\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11636_ _04746_ _04924_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__nor2_1
X_11567_ _05433_ _05467_ VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10518_ _04420_ _04421_ _04422_ _04423_ _00621_ VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__a221o_1
X_11498_ _05378_ _05398_ VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__xnor2_1
X_10449_ _04344_ _04354_ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__or2_1
X_12119_ _01578_ _04490_ VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07660_ _01720_ H\[3\]\[4\] _01629_ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__mux2_1
X_07591_ result_reg_mul\[2\] _01653_ _01561_ VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__o21ai_1
X_06611_ _00528_ _00631_ _00527_ _00634_ VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__or4_2
XFILLER_0_62_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06542_ _00568_ _00527_ _00665_ _00676_ _00603_ VGND VGND VPWR VPWR _00677_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_75_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09330_ _02687_ _02895_ VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09261_ R1\[0\] _00584_ VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__nand2_1
X_06473_ _00607_ VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__clkbuf_4
X_08212_ _00003_ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__clkbuf_4
X_09192_ _03102_ _02572_ _00586_ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08143_ H\[0\]\[13\] _01898_ _02074_ VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08074_ _01898_ H\[2\]\[13\] _02037_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07025_ _01127_ VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08976_ _02528_ H\[1\]\[3\] _02727_ VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07927_ CMD_setloop VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__clkbuf_4
X_07858_ _01906_ _01663_ _01907_ _01908_ VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_67_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06809_ _00931_ _00934_ _00732_ VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__mux2_1
X_07789_ _01841_ _01653_ _01842_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09528_ _01536_ _03423_ _03425_ _00549_ _03437_ VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__a311o_2
XFILLER_0_38_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09459_ _03225_ _03368_ VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__nor2_1
X_12470_ _06102_ _00647_ _06124_ _06171_ VGND VGND VPWR VPWR _06198_ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11421_ _05319_ _02486_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11352_ _05252_ _05253_ VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10303_ _04207_ _04209_ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11283_ _05183_ _05177_ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__nand2_1
X_13022_ clknet_leaf_28_clk _00465_ VGND VGND VPWR VPWR Qset\[3\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_10234_ _04117_ _04119_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__nand2_1
X_10165_ _04071_ _02573_ _00588_ VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__a21oi_1
X_10096_ _04001_ _04002_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__nand2_1
X_12806_ clknet_leaf_11_clk _00249_ VGND VGND VPWR VPWR result_reg_add\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10998_ _04096_ _03506_ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12737_ clknet_leaf_26_clk _00180_ VGND VGND VPWR VPWR H\[2\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12668_ clknet_leaf_42_clk _00118_ VGND VGND VPWR VPWR Oset\[2\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_11619_ _05415_ _05418_ _05417_ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12599_ clknet_leaf_39_clk _00049_ VGND VGND VPWR VPWR Qset\[1\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08830_ _02704_ _02743_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08761_ _02185_ _00583_ _02571_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__a21oi_1
X_07712_ net14 _01635_ VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__nor2_1
X_08692_ _02606_ VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__inv_2
X_07643_ _01702_ _01549_ _01703_ VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07574_ _01636_ _01549_ _01637_ VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__a21o_1
X_09313_ _03176_ _03080_ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__nand2_1
X_06525_ _00658_ _00659_ _00643_ VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06456_ _00590_ VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__inv_4
X_09244_ _02560_ _03151_ _03153_ _03154_ VGND VGND VPWR VPWR _03155_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_7_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09175_ _03085_ _02796_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06387_ _00520_ _00475_ _00522_ next_PC\[9\] _00478_ VGND VGND VPWR VPWR _00023_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08126_ _02080_ VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08057_ _02043_ VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07008_ _01118_ VGND VGND VPWR VPWR _00048_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput48 net48 VGND VGND VPWR VPWR data_out[0] sky130_fd_sc_hd__buf_1
Xoutput37 net37 VGND VGND VPWR VPWR data_W sky130_fd_sc_hd__buf_1
Xoutput59 net59 VGND VGND VPWR VPWR data_out[5] sky130_fd_sc_hd__buf_1
X_08959_ _00580_ _00671_ _02539_ VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__o21ai_2
X_11970_ _05811_ VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__inv_2
X_10921_ _04641_ _04636_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__nand2_1
X_10852_ _04754_ _04561_ _04564_ VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10783_ _02419_ _00584_ _03768_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12522_ net73 _06220_ _06221_ _06230_ VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_51_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_93_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12453_ _06267_ Him VGND VGND VPWR VPWR _06184_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12384_ _06126_ _02118_ VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11404_ _05304_ _05305_ _05175_ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__nand3_1
X_11335_ _05236_ _05065_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11266_ _05164_ _05165_ _05166_ _05167_ _00647_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__a221o_1
X_10217_ _04096_ _02785_ VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__nand2_1
X_13005_ clknet_leaf_35_clk _00448_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dfxtp_1
X_11197_ _05098_ _05099_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__nand2_1
X_10148_ _03152_ _04053_ _04054_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__o21ai_1
X_10079_ _03961_ _03985_ VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06310_ _06271_ _06261_ VGND VGND VPWR VPWR _06272_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07290_ Oset\[3\]\[6\] _01368_ _01250_ VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_42_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09931_ _02565_ Qset\[0\]\[9\] VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09862_ _02345_ _00584_ _03768_ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__a21o_1
X_08813_ _00007_ VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__buf_4
X_09793_ _03683_ _03699_ _03700_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__nand3_1
X_08744_ _02581_ Qset\[0\]\[1\] VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08675_ _00005_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__clkinv_4
X_07626_ _01584_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__clkbuf_4
X_07557_ _01611_ _01620_ _01621_ _01568_ VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06508_ _00642_ VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_33_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07488_ _01552_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__clkbuf_4
X_06439_ Him _00571_ _00573_ VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__nor3_4
X_09227_ _02545_ H\[1\]\[5\] VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__nand2_1
X_09158_ _02874_ H\[0\]\[7\] VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08109_ _01898_ H\[1\]\[13\] _02056_ VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09089_ _02989_ _02999_ _02540_ VGND VGND VPWR VPWR _03000_ sky130_fd_sc_hd__nand3_1
XFILLER_0_101_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11120_ _05021_ _05022_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11051_ _03652_ _04096_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__nand2_1
X_10002_ _03908_ _03859_ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11953_ _03819_ _00590_ VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11884_ _05735_ _05736_ VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__nand2_1
X_10904_ Oset\[3\]\[11\] _03792_ _03795_ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__a21oi_1
X_10835_ _04729_ _02409_ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_24_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10766_ H\[2\]\[11\] H\[3\]\[11\] _03760_ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__mux2_1
X_12505_ next_PC\[0\] _06218_ VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__or2_1
X_10697_ _04600_ _04601_ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__nand2_1
X_12436_ _06255_ _06113_ VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_10_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12367_ net22 net23 VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_74_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12298_ _06063_ _06064_ VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__nand2_1
X_11318_ _05218_ _05219_ VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__nand2_1
X_11249_ _04832_ H\[0\]\[13\] VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06790_ net15 _00600_ _00916_ VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08460_ _02311_ _02363_ _02140_ _02371_ _02381_ VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__o221ai_4
X_07411_ _01264_ _01035_ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__nand2_1
X_08391_ Qset\[0\]\[7\] VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__inv_2
X_07342_ _01412_ _01417_ _01214_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07273_ result_reg_not\[6\] _01351_ _01168_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09012_ _02539_ _02923_ _01153_ VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09914_ _02562_ Oset\[0\]\[8\] VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09845_ _03280_ _03751_ _00831_ VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__a21o_1
X_06988_ _01107_ VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__clkbuf_1
X_09776_ _03543_ _03551_ _03554_ VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__o21a_1
X_08727_ _01536_ _02628_ _02630_ _00548_ _02641_ VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_44_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _02572_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__buf_4
XFILLER_0_95_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07609_ _01603_ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_105_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08589_ _02491_ Qset\[1\]\[15\] _02444_ _02504_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__a211o_1
XFILLER_0_91_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10620_ _04448_ _04524_ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10551_ _04278_ _04276_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_24_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10482_ _04386_ _04385_ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12221_ result_reg_or\[11\] _05959_ _05857_ _06012_ VGND VGND VPWR VPWR _00367_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12152_ _05954_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__inv_2
X_12083_ _02944_ _05898_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__nand2_1
X_11103_ _05004_ _05005_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__nand2_1
X_11034_ _04935_ _04936_ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__nand2_1
X_12985_ clknet_leaf_7_clk _00428_ VGND VGND VPWR VPWR Him sky130_fd_sc_hd__dfxtp_1
X_11936_ _05782_ VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11867_ _05706_ _04444_ VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11798_ _05669_ VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__clkbuf_4
X_10818_ _04721_ _03746_ VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__nand2_1
X_10749_ _04650_ _04652_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12419_ _06155_ _06156_ _02116_ VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__a21oi_1
X_07960_ _06280_ im_reg\[6\] _01960_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__mux2_1
X_06911_ result_reg_set\[13\] VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_4_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
X_07891_ _01225_ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__inv_2
X_06842_ result_reg_sub\[10\] _00740_ _00966_ VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__o21ai_1
X_09630_ _03381_ _03403_ VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__nor2_1
X_06773_ result_reg_Lshift\[7\] VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__inv_2
X_09561_ _03467_ _03468_ _03469_ VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__nand3_1
X_08512_ _02328_ Qset\[3\]\[12\] _02347_ _02430_ VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__a211o_1
XFILLER_0_77_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09492_ _03400_ _03397_ _03398_ VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_92_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08443_ Oset\[2\]\[9\] VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08374_ Oset\[0\]\[6\] VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_98_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07325_ _00919_ _01275_ _01276_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__a21oi_1
X_07256_ _00841_ _00812_ _01173_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07187_ _01261_ VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__buf_2
XFILLER_0_14_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09828_ _03729_ _03732_ _03596_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_100_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09759_ _03608_ _03666_ VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12770_ clknet_leaf_26_clk _00213_ VGND VGND VPWR VPWR H\[0\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11721_ _05492_ _05620_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__nand2_1
X_11652_ _05532_ _05551_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__xor2_1
XFILLER_0_49_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10603_ _04318_ _04505_ _04313_ VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__nand3_1
XFILLER_0_91_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11583_ _05314_ _05311_ _05313_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_51_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10534_ _04439_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10465_ _04368_ _04370_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__or2_1
X_12204_ _03775_ _03824_ VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__nand2_1
X_10396_ _03773_ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_71_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12135_ _05907_ _04963_ _05147_ _05878_ VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_102_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12066_ _01578_ _02730_ VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11017_ _04918_ _04919_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__nand2_1
Xclkbuf_3_7__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12968_ clknet_leaf_7_clk _00411_ VGND VGND VPWR VPWR CMD_addition sky130_fd_sc_hd__dfxtp_2
XFILLER_0_87_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ clknet_leaf_15_clk _00342_ VGND VGND VPWR VPWR result_reg_and\[2\] sky130_fd_sc_hd__dfxtp_1
X_11919_ _03162_ VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07110_ _01183_ _01187_ _01192_ _01194_ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08090_ _02061_ VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07041_ _00904_ Qset\[2\]\[7\] _01129_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08992_ _02895_ VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07943_ _01973_ VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__clkbuf_1
X_07874_ net7 _01746_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__nor2_1
X_06825_ result_reg_Rshift\[9\] _00753_ _00950_ VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__o21ai_1
X_09613_ _03225_ _03223_ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__or2_1
X_06756_ result_reg_add\[7\] VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09544_ _03269_ _03270_ _03361_ VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__nand3_1
X_06687_ result_reg_and\[5\] _00562_ _00709_ VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__o21ai_1
X_09475_ _03184_ _03076_ VGND VGND VPWR VPWR _03385_ sky130_fd_sc_hd__nand2_1
X_08426_ _02327_ _02346_ _02347_ _02348_ VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_102_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08357_ _02260_ _02281_ _02250_ _02282_ VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__a211o_1
X_07308_ Oset\[3\]\[7\] _01385_ _01250_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__mux2_1
X_08288_ _02151_ Qset\[2\]\[3\] VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__nand2_1
X_07239_ _00786_ _01319_ _01181_ VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10250_ _04155_ _04031_ _04040_ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__nand3b_2
X_10181_ _04081_ _01155_ _04087_ _03066_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_6_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12822_ clknet_leaf_10_clk _00265_ VGND VGND VPWR VPWR result_reg_sub\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12753_ clknet_leaf_26_clk _00196_ VGND VGND VPWR VPWR H\[1\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11704_ _04855_ Qset\[2\]\[15\] VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__nand2_1
X_12684_ clknet_leaf_1_clk _00134_ VGND VGND VPWR VPWR LC\[8\] sky130_fd_sc_hd__dfxtp_1
X_11635_ _03233_ _05534_ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11566_ _05465_ _05466_ _03048_ VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__nand3_1
XFILLER_0_52_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10517_ Qset\[1\]\[9\] _03792_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__nand2_1
X_11497_ _05396_ _05397_ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__xor2_1
X_10448_ _04352_ _04353_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10379_ _04283_ Oset\[3\]\[9\] _03761_ _04284_ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__a211o_1
X_12118_ _01200_ _04483_ _04546_ VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__or3_1
X_12049_ _05844_ _01102_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07590_ _01548_ VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__buf_2
X_06610_ _00561_ VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__buf_2
X_06541_ _00628_ _00560_ _00552_ VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06472_ _00579_ _00605_ _00606_ VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__or3_2
X_09260_ _03163_ _01155_ _03170_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__nand3_1
X_08211_ Oset\[2\]\[0\] VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09191_ _02535_ _03098_ _03099_ _03101_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__a31o_2
X_08142_ _02088_ VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_31_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08073_ _02051_ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07024_ _00684_ _01126_ VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08975_ _02798_ _02234_ VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__nor2_1
X_07926_ R3\[0\] VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07857_ result_reg_mul\[14\] _01688_ _01667_ VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_67_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06808_ _00932_ _00933_ _00730_ VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__mux2_1
X_07788_ result_reg_mul\[11\] _01679_ _01656_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__o21ai_1
X_06739_ _00867_ _00615_ VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09527_ _01536_ _03436_ VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09458_ _03367_ VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__inv_2
X_09389_ _03298_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__inv_2
X_08409_ _02327_ H\[1\]\[7\] _02332_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__o21ai_1
X_11420_ _05319_ Oset\[3\]\[14\] _04303_ _05320_ VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11351_ _05251_ _05250_ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10302_ _04208_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__inv_2
X_11282_ _05177_ _05183_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__nor2_1
X_13021_ clknet_leaf_29_clk _00464_ VGND VGND VPWR VPWR Qset\[3\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_10233_ _04139_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10164_ _02560_ _04067_ _04068_ _04070_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__o31a_2
X_10095_ _04000_ _03997_ _03998_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_88_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12805_ clknet_leaf_11_clk _00248_ VGND VGND VPWR VPWR result_reg_add\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10997_ _04768_ _04765_ _04767_ VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12736_ clknet_leaf_33_clk _00179_ VGND VGND VPWR VPWR H\[2\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12667_ clknet_leaf_41_clk _00117_ VGND VGND VPWR VPWR Oset\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11618_ _05517_ _04896_ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__nand2_1
X_12598_ clknet_leaf_40_clk _00048_ VGND VGND VPWR VPWR Qset\[1\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_11549_ _05448_ _05438_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_77_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08760_ _02664_ _02673_ VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__nand2_1
X_07711_ _00881_ _01561_ VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__or2_1
X_08691_ _02605_ _01153_ VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__nand2_1
X_07642_ result_reg_mul\[4\] _01679_ _01561_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_0_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07573_ result_reg_mul\[1\] _01549_ _01561_ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__o21ai_1
X_09312_ _03222_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__inv_2
X_06524_ result_reg_Lshift\[0\] VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06455_ _00585_ _00589_ VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__nor2_4
X_09243_ _02567_ H\[3\]\[4\] _03135_ VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__a21oi_1
X_06386_ _06285_ _00521_ VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09174_ _03082_ _03084_ _00581_ VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__nand3_1
XFILLER_0_105_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_444 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08125_ H\[0\]\[4\] _01720_ _02075_ VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08056_ _01720_ H\[2\]\[4\] _02038_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput38 net38 VGND VGND VPWR VPWR data_address[0] sky130_fd_sc_hd__buf_1
X_07007_ _00927_ Qset\[1\]\[8\] _01109_ VGND VGND VPWR VPWR _01118_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput49 net49 VGND VGND VPWR VPWR data_out[10] sky130_fd_sc_hd__buf_1
X_08958_ _02866_ _02869_ _00581_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__nand3_1
X_07909_ _01950_ VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__clkbuf_1
X_08889_ _02522_ Oset\[0\]\[2\] VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__nand2_1
X_10920_ _04822_ _04823_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__nand2_2
X_10851_ _04561_ _04564_ _04754_ VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__a21o_1
X_10782_ _03770_ _04672_ _04678_ _04685_ VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12521_ _06219_ _00515_ VGND VGND VPWR VPWR _06230_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12452_ _06126_ _06182_ _04827_ _06183_ VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11403_ _00820_ _04974_ _02160_ _05299_ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__o211ai_1
X_12383_ _06267_ VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__buf_2
X_11334_ _03652_ _03110_ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__nand2_1
X_11265_ Oset\[1\]\[13\] _04857_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__nand2_1
X_10216_ _02949_ _04050_ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__nor2_1
X_13004_ clknet_leaf_36_clk _00447_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dfxtp_1
X_11196_ _05097_ _05092_ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__nand2_1
X_10147_ _03136_ Qset\[0\]\[14\] _02526_ VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10078_ _03984_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_12719_ clknet_leaf_36_clk _00162_ VGND VGND VPWR VPWR Oset\[1\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09930_ _03157_ Qset\[2\]\[9\] _02526_ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09861_ _02573_ VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__buf_4
X_08812_ _02561_ _02186_ _02725_ VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__o21ai_1
X_09792_ _03698_ _03684_ VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__nand2_1
X_08743_ _02655_ _00005_ _02656_ VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__nand3_1
XFILLER_0_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ _02581_ Qset\[0\]\[0\] VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__nand2_1
X_07625_ _01586_ result_reg_sub\[3\] VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07556_ _01571_ _00565_ _01540_ _01579_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__a211o_1
X_06507_ _00530_ _00592_ _00641_ VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09226_ _03136_ H\[0\]\[5\] VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__nand2_1
X_07487_ _01551_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__buf_4
XFILLER_0_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06438_ _00572_ VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__inv_2
X_09157_ _03065_ _03067_ VGND VGND VPWR VPWR _03068_ sky130_fd_sc_hd__nand2_1
X_06369_ _00507_ VGND VGND VPWR VPWR _00508_ sky130_fd_sc_hd__inv_2
X_08108_ _02070_ VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09088_ _02998_ _00581_ VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__nand2_1
X_08039_ Oset\[1\]\[13\] _01490_ _02018_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11050_ _04951_ _04952_ _03751_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__a21o_1
X_10001_ _03049_ _02738_ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__nor2_1
X_11952_ _03824_ _01158_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11883_ result_reg_mac\[14\] _05703_ _01149_ VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__o21a_1
X_10903_ Oset\[1\]\[11\] _03792_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__nand2_1
X_10834_ _04729_ Qset\[3\]\[11\] _04045_ _04737_ VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12504_ _06259_ VGND VGND VPWR VPWR _06221_ sky130_fd_sc_hd__clkbuf_4
X_10765_ _02423_ _04283_ _03764_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10696_ _04598_ _04528_ _04530_ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__nand3_1
XFILLER_0_42_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12435_ _01146_ _01554_ _06167_ _06160_ _06168_ VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12366_ _06097_ _02160_ _04827_ _06111_ VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__o211a_1
X_11317_ _04895_ _05158_ _05217_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12297_ _05766_ _03172_ _01959_ _02126_ _03175_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__o221a_1
X_11248_ _05142_ _05149_ _00585_ _02466_ VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__a2bb2o_1
X_11179_ _05062_ _05081_ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07410_ result_reg_and\[13\] _01207_ _01261_ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__o21a_1
X_08390_ _02248_ Qset\[3\]\[7\] _02254_ _02313_ VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__a211o_1
X_07341_ _01415_ _01193_ _01191_ _01416_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__a211o_1
XFILLER_0_73_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07272_ result_reg_Lshift\[6\] result_reg_Rshift\[6\] _01165_ VGND VGND VPWR VPWR
+ _01351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09011_ _02919_ _02922_ VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09913_ _02162_ _03819_ _02542_ VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09844_ _03047_ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__buf_4
X_06987_ _01106_ Qset\[0\]\[15\] _00686_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__mux2_1
X_09775_ _03562_ _03559_ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__nand2_1
X_08726_ Oreg3 _02635_ _00626_ _02640_ VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08657_ _02571_ VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__buf_6
X_07608_ _01670_ result_reg_mac\[2\] _01570_ VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ _02470_ _02503_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07539_ _01603_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10550_ _04318_ _04313_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_24_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10481_ _04367_ _04385_ _04386_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__nand3_1
X_09209_ _02798_ _02274_ VGND VGND VPWR VPWR _03120_ sky130_fd_sc_hd__nor2_1
X_12220_ _05937_ _06009_ _06010_ _06011_ _05957_ VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_102_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12151_ _00554_ _05666_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__nor2_1
X_12082_ _05888_ _02891_ VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__nor2_1
X_11102_ _04895_ _04924_ _05003_ VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__o21ai_1
X_11033_ _04934_ _04927_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__nand2_1
X_12984_ clknet_leaf_2_clk _00427_ VGND VGND VPWR VPWR Hreg3 sky130_fd_sc_hd__dfxtp_2
X_11935_ _00806_ _05774_ _05775_ _05781_ VGND VGND VPWR VPWR _05782_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11866_ _05724_ VGND VGND VPWR VPWR _00300_ sky130_fd_sc_hd__inv_2
X_11797_ result_reg_mul\[3\] _05670_ _05672_ _05676_ VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__o211a_1
X_10817_ _04719_ _04720_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__nand2_1
X_10748_ _03790_ _04651_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12418_ _06126_ CMD_store VGND VGND VPWR VPWR _06156_ sky130_fd_sc_hd__nand2_1
X_10679_ _04582_ _04576_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12349_ _01146_ VGND VGND VPWR VPWR _06097_ sky130_fd_sc_hd__buf_2
XFILLER_0_49_22 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06910_ net5 VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__inv_2
X_07890_ _01939_ VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__clkbuf_1
X_06841_ _00540_ _00959_ _00534_ VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06772_ result_reg_Rshift\[7\] VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__inv_2
X_09560_ _03421_ _03304_ VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__nand2_1
X_08511_ _02328_ _02429_ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__nor2_1
X_09491_ _03399_ _03400_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__nand2_1
X_08442_ _02328_ VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__buf_4
XFILLER_0_46_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08373_ _02261_ Oset\[3\]\[6\] _02254_ _02297_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__a211o_1
XFILLER_0_18_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07324_ _01254_ _01389_ _01394_ _01400_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__a31o_1
X_07255_ result_reg_not\[5\] _01334_ _01168_ VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07186_ result_reg_mul\[1\] _01263_ _01245_ _01269_ VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__a211o_1
XFILLER_0_41_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09827_ _03733_ _03734_ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__nand2_1
X_09758_ _03664_ _03665_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08709_ _00000_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__clkbuf_4
X_11720_ _05619_ VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__inv_2
X_09689_ _03444_ _03597_ VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__nor2_1
X_11651_ _05533_ _05550_ VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__xor2_1
XFILLER_0_36_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11582_ _05481_ _05482_ VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__nand2_1
X_10602_ _04455_ _04506_ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10533_ _04437_ _04435_ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10464_ _04369_ _04124_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__xor2_1
X_12203_ _03831_ _03767_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__nand2_1
X_10395_ _04283_ H\[0\]\[9\] VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_71_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12134_ result_reg_and\[12\] _05894_ _05936_ _05939_ _05940_ VGND VGND VPWR VPWR
+ _00352_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12065_ _05881_ _05882_ _02719_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__or3_1
X_11016_ _04917_ _04916_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12967_ clknet_leaf_6_clk _00410_ VGND VGND VPWR VPWR im_reg\[9\] sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_82_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12898_ clknet_leaf_14_clk _00341_ VGND VGND VPWR VPWR result_reg_and\[1\] sky130_fd_sc_hd__dfxtp_1
X_11918_ _05749_ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__buf_4
X_11849_ _05706_ _02986_ VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07040_ _01136_ VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08991_ _02618_ _02158_ _02897_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__a21oi_1
X_07942_ _01972_ LC\[2\] _01964_ VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__mux2_1
X_07873_ _01092_ _01560_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__or2_1
X_06824_ _00754_ _00949_ VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__nand2_1
X_09612_ _03519_ _03520_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09543_ _03447_ _03291_ _03446_ VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__a21oi_4
X_06755_ result_reg_sub\[7\] VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06686_ _00815_ _00745_ VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__or2_1
X_09474_ _03205_ _03383_ VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__nor2_1
X_08425_ H\[3\]\[8\] _02327_ VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_102_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08356_ H\[1\]\[5\] _02230_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__nor2_1
X_07307_ _01161_ _01371_ _01383_ _01384_ VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__a22o_4
XFILLER_0_18_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08287_ _02215_ VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__clkbuf_1
X_07238_ _00787_ _01318_ _01176_ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__mux2_1
X_07169_ result_reg_not\[1\] _01252_ _01168_ VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__mux2_1
X_10180_ _04086_ _02552_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_6_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12821_ clknet_leaf_11_clk _00264_ VGND VGND VPWR VPWR result_reg_sub\[4\] sky130_fd_sc_hd__dfxtp_1
X_12752_ clknet_leaf_33_clk _00195_ VGND VGND VPWR VPWR H\[1\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_11703_ _03795_ _05600_ _05601_ _05602_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__a2bb2o_1
X_12683_ clknet_leaf_1_clk _00133_ VGND VGND VPWR VPWR LC\[7\] sky130_fd_sc_hd__dfxtp_1
X_11634_ _05341_ _03859_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11565_ _05463_ _05205_ _05201_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__nand3_1
XFILLER_0_4_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11496_ _05279_ _05272_ VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__nand2_1
X_10516_ _04414_ Qset\[0\]\[9\] _03798_ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__a21oi_1
X_10447_ _04351_ _04346_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__nand2_1
X_10378_ _04283_ _02365_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__nor2_1
X_12117_ _01407_ _05873_ _02115_ _05926_ VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__a211oi_1
X_12048_ result_reg_Rshift\[14\] _05848_ _05857_ _05868_ VGND VGND VPWR VPWR _00338_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06540_ _00669_ _00665_ _00674_ VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__o21a_1
X_06471_ _00530_ _00528_ VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08210_ _02127_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__buf_6
XFILLER_0_28_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09190_ _02787_ H\[2\]\[6\] _03100_ VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__a21oi_1
X_08141_ H\[0\]\[12\] _01879_ _02074_ VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08072_ _01879_ H\[2\]\[12\] _02037_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07023_ _00675_ _00677_ VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__or2b_1
XFILLER_0_11_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08974_ _02883_ _02885_ VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07925_ _01958_ VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__clkbuf_1
X_07856_ _01579_ result_reg_sub\[14\] VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_3_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06807_ result_reg_add\[9\] VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__inv_2
X_07787_ _00991_ _00982_ _01544_ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06738_ _00860_ _00866_ _00732_ VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09526_ _03430_ _03435_ _00646_ VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__mux2_1
X_09457_ _03176_ _03052_ _03220_ VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06669_ _00797_ _00743_ _00798_ _00799_ VGND VGND VPWR VPWR _00800_ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08408_ _02319_ H\[0\]\[7\] _02254_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__o21a_1
X_09388_ _03289_ _03297_ VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08339_ _02265_ net58 _02170_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__mux2_1
X_11350_ _05250_ _05251_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10301_ _03651_ _03304_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13020_ clknet_leaf_35_clk _00463_ VGND VGND VPWR VPWR Qset\[3\]\[11\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_5_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11281_ _05181_ _05182_ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__xnor2_1
X_10232_ _04137_ _04120_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10163_ _02490_ _03157_ _03135_ _04069_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__a211o_1
X_10094_ _03999_ _04000_ VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12804_ clknet_leaf_11_clk _00247_ VGND VGND VPWR VPWR result_reg_add\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10996_ _04896_ _03079_ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__nand2_2
X_12735_ clknet_leaf_33_clk _00178_ VGND VGND VPWR VPWR H\[2\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12666_ clknet_leaf_44_clk _00116_ VGND VGND VPWR VPWR Oset\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11617_ _05516_ _01554_ _02519_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__a21bo_2
X_12597_ clknet_leaf_43_clk _00047_ VGND VGND VPWR VPWR Qset\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11548_ _05438_ _05448_ VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__or2_1
X_11479_ _04281_ _05379_ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_90_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07710_ _01766_ _01549_ _01767_ VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__a21o_1
X_08690_ _02601_ _02604_ _02551_ VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__nand3_1
X_07641_ _00788_ _00789_ _01545_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_69_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07572_ _00702_ _00703_ _01545_ VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06523_ result_reg_Rshift\[0\] VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__inv_2
X_09311_ _03178_ _03221_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__xor2_1
XFILLER_0_75_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06454_ _00588_ VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__buf_4
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09242_ _03152_ H\[2\]\[4\] VGND VGND VPWR VPWR _03153_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06385_ next_PC\[9\] _00516_ VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__xor2_1
X_09173_ _02544_ Qset\[3\]\[6\] _02800_ _03083_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__a211o_1
X_08124_ _02079_ VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_78_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08055_ _02042_ VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput39 net39 VGND VGND VPWR VPWR data_address[1] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_8_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07006_ _01117_ VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08957_ _02867_ _02800_ _02868_ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_87_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07908_ Oset\[2\]\[7\] _01385_ _01942_ VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__mux2_1
X_08888_ _02799_ _02800_ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__nand2_1
X_07839_ _01571_ _00551_ _01042_ _01588_ VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_98_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10850_ _04725_ _04753_ VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__xor2_1
XFILLER_0_85_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09509_ _03383_ _00556_ VGND VGND VPWR VPWR _03419_ sky130_fd_sc_hd__nand2_1
X_10781_ _00584_ _04684_ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__or2_1
X_12520_ net72 _06220_ _06221_ _06229_ VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12451_ _06126_ _00626_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11402_ _05300_ _00832_ VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_90 _01775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12382_ _06114_ net23 _06116_ _06124_ VGND VGND VPWR VPWR _06125_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11333_ _03652_ _03076_ VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__nand2_1
X_11264_ _04415_ Oset\[0\]\[13\] _04862_ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__a21oi_1
X_10215_ _04098_ _04051_ _04121_ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__a21oi_1
X_13003_ clknet_leaf_38_clk _00446_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dfxtp_1
X_11195_ _05092_ _05097_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__or2_1
X_10146_ Qset\[1\]\[14\] VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10077_ _03982_ _03983_ VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10979_ _04881_ Oset\[1\]\[12\] VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12718_ clknet_leaf_40_clk _00161_ VGND VGND VPWR VPWR Oset\[1\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_12649_ clknet_leaf_41_clk _00099_ VGND VGND VPWR VPWR H\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09860_ _03763_ _03766_ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__nand2_2
XFILLER_0_0_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08811_ _02527_ H\[3\]\[1\] VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__nand2_1
X_09791_ _03684_ _03698_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__or2_1
X_08742_ _02585_ Qset\[3\]\[1\] VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08673_ _02583_ _02584_ _02587_ VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__nand3_1
X_07624_ _01581_ result_reg_add\[3\] VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_49_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07555_ _01583_ _01573_ _01588_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__or3b_1
XFILLER_0_48_334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06506_ _00638_ shift.left _00637_ VGND VGND VPWR VPWR _00641_ sky130_fd_sc_hd__and3_2
XFILLER_0_48_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07486_ _00586_ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__inv_2
X_09225_ _02787_ VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__buf_4
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06437_ Qreg2 _00525_ VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__nor2_2
XFILLER_0_33_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09156_ _03066_ VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06368_ _00506_ _00501_ VGND VGND VPWR VPWR _00507_ sky130_fd_sc_hd__or2_1
X_08107_ _01879_ H\[1\]\[12\] _02056_ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06299_ current_state\[5\] VGND VGND VPWR VPWR _06264_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09087_ _02994_ _02997_ VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__nand2_1
X_08038_ _02032_ VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10000_ _03906_ VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_95_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09989_ _03894_ _03895_ VGND VGND VPWR VPWR _03896_ sky130_fd_sc_hd__nand2_1
X_11951_ result_reg_Lshift\[6\] _05743_ _05672_ _05795_ VGND VGND VPWR VPWR _00314_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11882_ _05485_ _05486_ _05703_ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__nand3_1
X_10902_ _04414_ Oset\[0\]\[11\] VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10833_ _04729_ _02406_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10764_ _04302_ _03861_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12503_ _06219_ VGND VGND VPWR VPWR _06220_ sky130_fd_sc_hd__clkbuf_4
X_10695_ _04531_ _04599_ VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12434_ _06165_ _06149_ _06124_ VGND VGND VPWR VPWR _06168_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12365_ _06110_ _06097_ VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11316_ _04895_ _05158_ _05217_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_74_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12296_ _06058_ VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__buf_2
X_11247_ _05147_ _00582_ _03781_ _05148_ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__a211oi_1
X_11178_ _05077_ _05080_ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__nand2_1
X_10129_ _04006_ VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07340_ net16 _01186_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07271_ _01350_ VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__clkbuf_1
X_09010_ _02920_ _02590_ _02921_ VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__nand3_1
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09912_ _03815_ _03816_ _03817_ _03818_ VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__o22a_2
X_09843_ _03739_ _03749_ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__nand2_1
X_06986_ _01100_ _01105_ VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__nand2_1
X_09774_ _03676_ _03681_ _03274_ VGND VGND VPWR VPWR _03682_ sky130_fd_sc_hd__nand3_1
X_08725_ _02637_ _02639_ _00646_ VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__a21o_1
X_08656_ _02555_ VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__inv_6
X_07607_ _01594_ _01660_ _01669_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__o21ai_1
X_08587_ Qset\[0\]\[15\] VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_105_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07538_ _01602_ _01556_ VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_105_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07469_ _01534_ _01532_ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10480_ _04384_ _04383_ VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__or2_1
X_09208_ _03118_ VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09139_ _03049_ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__inv_6
XFILLER_0_32_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12150_ result_reg_and\[15\] _05894_ _05950_ _05953_ _05940_ VGND VGND VPWR VPWR
+ _00355_ sky130_fd_sc_hd__o221a_1
X_11101_ _04895_ _04924_ _05003_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__or3_1
XFILLER_0_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12081_ _05892_ _02933_ _05760_ VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11032_ _04927_ _04934_ VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12983_ clknet_leaf_7_clk _00426_ VGND VGND VPWR VPWR Hreg2 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_99_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11934_ _05774_ _05780_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_43_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _04257_ _05703_ _05710_ _05723_ VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11796_ _02957_ _05670_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__nand2_1
X_10816_ _04717_ _04526_ _04645_ VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__nand3_1
XFILLER_0_82_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10747_ _03897_ _02904_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10678_ _04576_ _04582_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12417_ _06266_ _06154_ _06151_ VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__or3_1
XFILLER_0_23_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12348_ _06096_ VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12279_ _06032_ _01101_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06840_ result_reg_or\[10\] VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06771_ result_reg_not\[7\] VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__inv_2
X_08510_ Qset\[2\]\[12\] VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__inv_2
X_09490_ _03350_ _03206_ VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08441_ _02359_ _02362_ VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__nand2_2
XFILLER_0_105_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08372_ _02248_ _02296_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_98_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07323_ _01398_ _01192_ _01399_ _01220_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__a31o_1
X_07254_ result_reg_Lshift\[5\] result_reg_Rshift\[5\] _01165_ VGND VGND VPWR VPWR
+ _01334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07185_ result_reg_add\[1\] _01264_ _01266_ _01268_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09826_ _03596_ VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__inv_2
X_06969_ _01085_ _00562_ _01087_ _01088_ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__a31o_1
X_09757_ _03662_ _03655_ _03658_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_57_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _02160_ _02622_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__xor2_4
XTAP_TAPCELL_ROW_29_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _03592_ _03596_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__nand2_1
X_08639_ _02543_ _02553_ VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11650_ _05547_ _05549_ VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__xor2_1
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11581_ _05306_ _05476_ _05479_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__nand3b_2
X_10601_ _04505_ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10532_ _04435_ _04437_ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10463_ _04074_ _02963_ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12202_ _05960_ _05996_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_23_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10394_ H\[2\]\[9\] H\[3\]\[9\] _04282_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12133_ _05682_ VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12064_ _02667_ _02670_ VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__nand2_1
X_11015_ _04916_ _04917_ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_32_Left_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12966_ clknet_leaf_6_clk _00409_ VGND VGND VPWR VPWR im_reg\[8\] sky130_fd_sc_hd__dfxtp_4
X_11917_ _00591_ _05754_ VGND VGND VPWR VPWR _05765_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_82_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ clknet_leaf_16_clk _00340_ VGND VGND VPWR VPWR result_reg_and\[0\] sky130_fd_sc_hd__dfxtp_1
X_11848_ _05712_ VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11779_ _05621_ _05622_ _05655_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__nand3_1
XFILLER_0_42_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_41_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_8 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08990_ _02896_ _02900_ _02901_ VGND VGND VPWR VPWR _02902_ sky130_fd_sc_hd__nand3_1
XFILLER_0_76_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07941_ _01971_ R2\[0\] _01960_ VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07872_ _01920_ _01653_ _01921_ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__a21o_1
X_06823_ result_reg_Lshift\[9\] VGND VGND VPWR VPWR _00949_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_50_Left_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09611_ _03518_ _03453_ _03456_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__nand3b_1
X_06754_ result_reg_mul\[7\] VGND VGND VPWR VPWR _00882_ sky130_fd_sc_hd__inv_2
X_09542_ _03451_ VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06685_ result_reg_mul\[5\] VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__inv_2
X_09473_ _03145_ VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__inv_2
X_08424_ _02254_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_102_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08355_ H\[0\]\[5\] VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__inv_2
X_07306_ _00880_ _01275_ _01276_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__a21oi_1
X_08286_ _02214_ net56 _02170_ VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07237_ _00788_ _00789_ _01173_ VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__mux2_1
X_07168_ result_reg_Lshift\[1\] result_reg_Rshift\[1\] _01165_ VGND VGND VPWR VPWR
+ _01252_ sky130_fd_sc_hd__mux2_1
X_07099_ _00698_ _00653_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__nor2_1
X_09809_ _03022_ Oset\[2\]\[7\] VGND VGND VPWR VPWR _03717_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_6_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12820_ clknet_leaf_11_clk _00263_ VGND VGND VPWR VPWR result_reg_sub\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12751_ clknet_leaf_33_clk _00194_ VGND VGND VPWR VPWR H\[1\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_11702_ _04415_ Oset\[0\]\[15\] _03798_ VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__a21oi_1
X_12682_ clknet_leaf_1_clk _00132_ VGND VGND VPWR VPWR LC\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11633_ _05436_ _05454_ _05457_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__o21ai_1
X_11564_ _05434_ _05464_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11495_ _05394_ _05395_ VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__nand2_1
X_10515_ _04414_ Qset\[2\]\[9\] VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__nand2_1
X_10446_ _04346_ _04351_ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10377_ _04282_ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__buf_6
X_12116_ _05923_ _05924_ _05925_ _05871_ VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__and4_1
X_12047_ _05839_ _05851_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12949_ clknet_leaf_15_clk _00392_ VGND VGND VPWR VPWR result_reg_set\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06470_ _00550_ _00592_ VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__nand2_1
XANTENNA_180 _02526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08140_ _02087_ VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08071_ _02050_ VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__clkbuf_1
X_07022_ _01125_ VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08973_ _02884_ VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__inv_2
X_07924_ Oset\[2\]\[15\] _01525_ _01941_ VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07855_ _01580_ result_reg_add\[14\] VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_3_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06806_ result_reg_sub\[9\] VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07786_ _01840_ VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_39_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06737_ _00865_ _00857_ _00730_ VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09525_ _03431_ _03432_ _02837_ _03433_ _03434_ VGND VGND VPWR VPWR _03435_ sky130_fd_sc_hd__a32o_1
X_06668_ result_reg_and\[4\] _00561_ _00552_ VGND VGND VPWR VPWR _00799_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_66_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09456_ _03362_ _03365_ VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__nand2_1
X_08407_ _02327_ H\[3\]\[7\] _02330_ VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06599_ _00613_ VGND VGND VPWR VPWR _00732_ sky130_fd_sc_hd__clkbuf_4
X_09387_ _03279_ _03296_ VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08338_ _02126_ _02247_ _02140_ _02257_ _02264_ VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_34_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08269_ _02128_ Qset\[0\]\[2\] VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11280_ _04854_ _03079_ _03859_ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__and3_1
X_10300_ _04203_ _04206_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__nor2_1
X_10231_ _04120_ _04137_ VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__nor2_1
X_10162_ _03157_ H\[2\]\[14\] VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10093_ _03897_ _03899_ _03685_ VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12803_ clknet_leaf_11_clk _00246_ VGND VGND VPWR VPWR result_reg_add\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_54_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_8
X_12734_ clknet_leaf_40_clk _00177_ VGND VGND VPWR VPWR H\[2\]\[9\] sky130_fd_sc_hd__dfxtp_2
X_10995_ _04772_ _04763_ _04771_ VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12665_ clknet_leaf_45_clk _00115_ VGND VGND VPWR VPWR Oset\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11616_ _05509_ _05515_ _03768_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__mux2_1
X_12596_ clknet_leaf_43_clk _00046_ VGND VGND VPWR VPWR Qset\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11547_ _05446_ _05447_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11478_ _05341_ VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_90_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10429_ _04333_ _04334_ _04246_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07640_ _01701_ VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__clkbuf_1
X_07571_ _01559_ VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_88_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06522_ _00656_ VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_45_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_8
X_09310_ _03220_ _03111_ _03180_ VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__o21ai_1
X_09241_ _02523_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__buf_4
X_06453_ _00587_ VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__clkbuf_4
X_06384_ im_reg\[9\] _06285_ VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__or2_1
X_09172_ _02528_ _02289_ VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08123_ H\[0\]\[3\] _01700_ _02075_ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08054_ _01700_ H\[2\]\[3\] _02038_ VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07005_ _00904_ Qset\[1\]\[7\] _01109_ VGND VGND VPWR VPWR _01117_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08956_ _02528_ Qset\[1\]\[3\] VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__nand2_1
X_07907_ _01949_ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__clkbuf_1
X_08887_ _02534_ VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__buf_6
X_07838_ _01887_ _01663_ _01888_ _01889_ VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__a31o_1
X_07769_ _00956_ _01682_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__or2_1
X_09508_ _03416_ _00623_ _03417_ VGND VGND VPWR VPWR _03418_ sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_36_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_8
X_10780_ _02540_ _04683_ VGND VGND VPWR VPWR _04684_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09439_ _03348_ _02286_ VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__nand2_2
X_12450_ _06130_ _06181_ VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__nor2_1
X_11401_ _05175_ _05301_ _05302_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__nand3b_1
XANTENNA_80 _01690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 _01788_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12381_ _06123_ current_state\[2\] VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__nand2_2
X_11332_ _03383_ _05063_ VGND VGND VPWR VPWR _05234_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11263_ _04415_ Oset\[2\]\[13\] VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__nand2_1
X_11194_ _04650_ _05093_ _05096_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__o21a_1
X_13002_ clknet_leaf_38_clk _00445_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dfxtp_1
X_10214_ _04075_ _04097_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__nor2_1
X_10145_ _04051_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__inv_2
X_10076_ _03976_ _03978_ _03980_ VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__nand3_2
XFILLER_0_85_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10978_ _04729_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__buf_4
XFILLER_0_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12717_ clknet_leaf_41_clk _00160_ VGND VGND VPWR VPWR Oset\[1\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_12648_ clknet_leaf_32_clk _00098_ VGND VGND VPWR VPWR H\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12579_ clknet_leaf_45_clk _00029_ VGND VGND VPWR VPWR Qset\[0\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08810_ _02721_ _02723_ VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09790_ _03686_ _03697_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__xor2_1
X_08741_ _02581_ Qset\[2\]\[1\] VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__nand2_1
X_08672_ _02586_ Qset\[3\]\[0\] VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__nand2_1
X_07623_ _01681_ _01635_ _01683_ _01684_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_49_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07554_ _01616_ _01618_ _00669_ _01606_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__o2bb2a_1
X_07485_ _01546_ _01549_ VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06505_ _00637_ _00639_ VGND VGND VPWR VPWR _00640_ sky130_fd_sc_hd__nor2_2
XFILLER_0_48_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06436_ _00570_ Qim VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__nand2_1
X_09224_ _02800_ VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__buf_4
XFILLER_0_33_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09155_ _01154_ _01990_ _02555_ VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_44_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06367_ next_PC\[6\] VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06298_ current_state\[0\] VGND VGND VPWR VPWR _06263_ sky130_fd_sc_hd__inv_2
X_09086_ _02995_ _02591_ _02996_ VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__nand3_1
X_08106_ _02069_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__clkbuf_1
X_08037_ Oset\[1\]\[12\] _01473_ _02018_ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09988_ _03892_ _03883_ _03884_ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__nand3_1
X_08939_ _00621_ _02846_ _02851_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__a21oi_1
X_11950_ _05794_ _05771_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__nand2_1
X_10901_ _04801_ _04802_ _03795_ _04803_ _04804_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__a32o_1
X_11881_ _05734_ VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10832_ _04735_ _03781_ _00585_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10763_ _04665_ _04666_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12502_ _06218_ VGND VGND VPWR VPWR _06219_ sky130_fd_sc_hd__inv_2
X_10694_ _04598_ VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12433_ _06164_ _06112_ VGND VGND VPWR VPWR _06167_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_10_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12364_ _06100_ _06099_ _06105_ _06106_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__a211o_1
X_11315_ _05215_ _05216_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12295_ _06061_ _06062_ _02116_ VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__a21oi_1
X_11246_ _02458_ _02163_ VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11177_ _04025_ _05079_ _05076_ VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__o21ai_1
X_10128_ _03960_ _04009_ _03985_ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__nand3b_1
X_10059_ _03965_ _03928_ VGND VGND VPWR VPWR _03966_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07270_ Oset\[3\]\[5\] _01349_ _01250_ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_7_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
X_09911_ Qset\[1\]\[8\] _03136_ _03135_ VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09842_ _03732_ _03734_ _03743_ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__a21oi_1
X_09773_ _03677_ _03680_ VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__nand2_1
X_06985_ _01101_ _00654_ _00656_ _01104_ _00665_ VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__a221o_1
X_08724_ Oset\[1\]\[0\] _02624_ _00001_ _02638_ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__a211o_1
XFILLER_0_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08655_ _02560_ _02564_ _02566_ _02569_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__o31ai_2
X_07606_ _00738_ _01574_ _01665_ _01668_ _01569_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08586_ _02491_ Qset\[3\]\[15\] _02374_ _02501_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_105_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07537_ _00641_ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_105_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07468_ R1\[1\] net30 current_state\[2\] VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__mux2_1
X_07399_ _01006_ _01275_ _01160_ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__a21oi_1
X_06419_ _00546_ VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09207_ _02544_ Oset\[1\]\[5\] VGND VGND VPWR VPWR _03118_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09138_ shift.H _02571_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__nor2_4
X_09069_ _02962_ _02980_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__nand2_1
X_11100_ _05001_ _05002_ VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__or2b_1
X_12080_ _05895_ _05894_ VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__nand2_1
X_11031_ _04932_ _04933_ VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__nand2_1
X_12982_ clknet_leaf_3_clk _00425_ VGND VGND VPWR VPWR shift.H sky130_fd_sc_hd__dfxtp_2
X_11933_ _05762_ _05776_ _02118_ _05779_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__o22ai_2
X_11864_ result_reg_mac\[8\] _05702_ VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_43_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10815_ _04646_ _04718_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11795_ result_reg_mul\[2\] _05670_ _05672_ _05675_ VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10746_ _04308_ _04460_ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10677_ _04577_ _04581_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_23_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12416_ _06104_ _06122_ _06253_ VGND VGND VPWR VPWR _06154_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12347_ _06095_ _01532_ VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12278_ _06039_ _05833_ _06044_ _06050_ VGND VGND VPWR VPWR _00386_ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11229_ _04876_ _05131_ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06770_ _00880_ _00725_ _00897_ VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08440_ _02356_ Qset\[1\]\[9\] _02329_ _02361_ VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__a211o_1
XFILLER_0_58_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08371_ Oset\[2\]\[6\] VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__inv_2
X_07322_ result_reg_or\[8\] _01199_ VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07253_ _01333_ VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07184_ _01267_ _00702_ VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09825_ _03729_ _03732_ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__nand2_1
X_06968_ result_reg_and\[15\] _00562_ _00709_ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__o21ai_1
X_09756_ _03659_ _03663_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_57_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _03593_ _03594_ _03595_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__nand3_1
X_08707_ _00622_ _02578_ _02621_ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__o21ai_4
X_06899_ _00739_ _01013_ _01015_ _01020_ _01021_ VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__a32o_1
X_08638_ _02550_ _02552_ VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08569_ Oset\[0\]\[14\] VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__inv_2
X_11580_ _05480_ _05306_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__nand2_1
X_10600_ _04502_ _04504_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10531_ _03756_ _03813_ _04436_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12201_ _03780_ _03819_ _05907_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10462_ _03205_ _04050_ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10393_ _01156_ _02371_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12132_ _05937_ _04886_ _04842_ _05938_ _04836_ VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__a32o_1
X_12063_ _01200_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11014_ _04762_ _04774_ _04776_ VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12965_ clknet_leaf_6_clk _00408_ VGND VGND VPWR VPWR im_reg\[7\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_35_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11916_ result_reg_Lshift\[2\] _05743_ _05672_ _05764_ VGND VGND VPWR VPWR _00310_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12896_ clknet_leaf_21_clk _00339_ VGND VGND VPWR VPWR result_reg_Rshift\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_82_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ _00724_ _05707_ _05710_ _05711_ VGND VGND VPWR VPWR _05712_ sky130_fd_sc_hd__a211o_1
XFILLER_0_74_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11778_ _05662_ VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10729_ _04631_ _04633_ VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07940_ _06274_ _01970_ VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__nand2_1
X_07871_ result_reg_mul\[15\] _01548_ _01656_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__o21ai_1
X_06822_ result_reg_not\[9\] VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__inv_2
X_09610_ _03457_ _03518_ VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__nand2_1
X_09541_ _00812_ _02654_ _02753_ _03450_ VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__a211o_1
X_06753_ result_reg_set\[7\] VGND VGND VPWR VPWR _00881_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06684_ result_reg_sub\[5\] _00541_ _00813_ VGND VGND VPWR VPWR _00814_ sky130_fd_sc_hd__o21ai_1
X_09472_ _03381_ VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08423_ H\[2\]\[8\] VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08354_ _02276_ _02279_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__nand2_1
X_07305_ _01254_ _01372_ _01376_ _01382_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__a31o_1
XFILLER_0_73_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08285_ _02126_ _02201_ _02140_ _02206_ _02213_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_33_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07236_ result_reg_not\[4\] _01316_ _01168_ VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07167_ _01251_ VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07098_ _01170_ _01178_ _01182_ VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__mux2_1
X_09808_ Oset\[3\]\[7\] _03033_ _03026_ VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_6_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09739_ _02991_ _03644_ _03645_ _03646_ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__o2bb2a_1
X_12750_ clknet_leaf_40_clk _00193_ VGND VGND VPWR VPWR H\[1\]\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_96_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11701_ Oset\[1\]\[15\] _04857_ VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__nand2_1
X_12681_ clknet_leaf_1_clk _00131_ VGND VGND VPWR VPWR LC\[5\] sky130_fd_sc_hd__dfxtp_1
X_11632_ _05465_ _05462_ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11563_ _05463_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11494_ _05391_ _05393_ _05392_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__nand3_1
X_10514_ Qset\[3\]\[9\] _03791_ _03794_ VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__a21oi_1
X_10445_ _04013_ _04347_ _04350_ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12115_ _00525_ _03840_ _04294_ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__or3_1
X_10376_ _03498_ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__buf_6
XFILLER_0_20_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12046_ result_reg_Rshift\[13\] _05848_ _05857_ _05867_ VGND VGND VPWR VPWR _00337_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12948_ clknet_leaf_14_clk _00391_ VGND VGND VPWR VPWR result_reg_set\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12879_ clknet_leaf_24_clk _00322_ VGND VGND VPWR VPWR result_reg_Lshift\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_170 _01332_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_181 _02526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08070_ _01859_ H\[2\]\[11\] _02037_ VGND VGND VPWR VPWR _02050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07021_ _01106_ Qset\[1\]\[15\] _01108_ VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08972_ _01153_ _00671_ _02555_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__o21ai_1
X_07923_ _01957_ VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__clkbuf_1
X_07854_ _01902_ _01658_ _01903_ _01904_ VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06805_ result_reg_mul\[9\] VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_3_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07785_ _01839_ H\[3\]\[10\] _01628_ VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06736_ result_reg_sub\[6\] VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09524_ _03021_ Qset\[2\]\[5\] VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__nand2_1
X_06667_ _00787_ _00745_ VGND VGND VPWR VPWR _00798_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09455_ _03363_ _03364_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__nand2_1
X_08406_ _02328_ H\[2\]\[7\] _02329_ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__o21a_1
X_06598_ _00728_ _00729_ _00730_ VGND VGND VPWR VPWR _00731_ sky130_fd_sc_hd__mux2_1
X_09386_ _00536_ _03280_ VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08337_ _02259_ _02263_ _01552_ VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__a21o_2
XFILLER_0_34_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08268_ _02195_ _00003_ _02196_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__nand3_1
XFILLER_0_104_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07219_ result_reg_add\[3\] _01267_ VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__nor2_1
X_10230_ _04135_ _04136_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__nand2_1
X_08199_ _02129_ Qset\[2\]\[0\] VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__nand2_1
X_10161_ H\[1\]\[14\] _03152_ VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__nor2_1
X_10092_ _03997_ _03998_ VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__nand2_1
X_12802_ clknet_leaf_9_clk _00245_ VGND VGND VPWR VPWR result_reg_add\[1\] sky130_fd_sc_hd__dfxtp_1
X_10994_ _04786_ _04780_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12733_ clknet_leaf_40_clk _00176_ VGND VGND VPWR VPWR H\[2\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12664_ clknet_leaf_43_clk _00114_ VGND VGND VPWR VPWR Oset\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_11615_ _04835_ _05510_ _05512_ _05514_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__o31a_1
X_12595_ clknet_leaf_45_clk _00045_ VGND VGND VPWR VPWR Qset\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11546_ _05445_ _05439_ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11477_ _05376_ _05377_ VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10428_ _04325_ _04327_ _04331_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__nand3_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10359_ _03651_ _03614_ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__nand2_2
X_12029_ _05794_ _05851_ VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07570_ _01633_ _00689_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_64_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06521_ _00636_ _00633_ VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__nand2_4
X_09240_ H\[0\]\[4\] H\[1\]\[4\] _02562_ VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06452_ _00586_ VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__buf_6
X_06383_ _00518_ _00475_ _00519_ next_PC\[8\] _00478_ VGND VGND VPWR VPWR _00022_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09171_ _02544_ Qset\[1\]\[6\] _02727_ _03081_ VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__a211o_1
XFILLER_0_7_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08122_ _02078_ VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08053_ _02041_ VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__clkbuf_1
X_07004_ _01116_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08955_ _02522_ Qset\[0\]\[3\] VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__nand2_1
X_07906_ Oset\[2\]\[6\] _01368_ _01942_ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__mux2_1
X_08886_ _02798_ Oset\[1\]\[2\] VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07837_ result_reg_mul\[13\] _01688_ _01667_ VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__o21ai_1
X_07768_ _01821_ _01653_ _01822_ VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__a21o_1
X_06719_ result_reg_not\[5\] VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09507_ _03407_ _03410_ _03233_ VGND VGND VPWR VPWR _03417_ sky130_fd_sc_hd__nand3_1
X_07699_ _01716_ _00874_ VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09438_ _03340_ _03347_ VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__nand2_2
XFILLER_0_93_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09369_ _00620_ _00523_ _00582_ VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12380_ net25 _06122_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__nor2_2
XFILLER_0_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11400_ _04830_ _04974_ _00832_ _05299_ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__o211ai_1
XANTENNA_81 _01711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_92 _01792_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_70 _01467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11331_ _05070_ _05066_ VGND VGND VPWR VPWR _05233_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11262_ Oset\[3\]\[13\] _04857_ _03795_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__a21oi_1
X_10213_ _04117_ _04118_ _04119_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__a21boi_1
X_13001_ clknet_leaf_39_clk _00444_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dfxtp_1
X_11193_ _05094_ _05095_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__nand2_1
X_10144_ _03115_ _04050_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10075_ _03979_ _03981_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10977_ _04879_ VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12716_ clknet_leaf_41_clk _00159_ VGND VGND VPWR VPWR Oset\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_550 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12647_ clknet_leaf_46_clk _00097_ VGND VGND VPWR VPWR H\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12578_ clknet_leaf_48_clk _00028_ VGND VGND VPWR VPWR Qset\[0\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_11529_ _05428_ _05429_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08740_ _02653_ VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__clkbuf_4
X_08671_ _02585_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__buf_6
X_07622_ net10 _01658_ VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07553_ R2\[1\] _01593_ _01540_ _01617_ VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__a211o_1
X_07484_ _01548_ VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__buf_2
X_06504_ _00638_ VGND VGND VPWR VPWR _00639_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06435_ Oim VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__inv_2
X_09223_ _03130_ _03133_ VGND VGND VPWR VPWR _03134_ sky130_fd_sc_hd__nand2_1
X_09154_ _03058_ _01154_ _03064_ VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__nand3_1
XFILLER_0_44_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06366_ im_reg\[6\] _06285_ VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__or2_1
X_08105_ _01859_ H\[1\]\[11\] _02056_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__mux2_1
X_06297_ _06262_ VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__inv_2
X_09085_ _02992_ Qset\[1\]\[4\] VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__nand2_1
X_08036_ _02031_ VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09987_ _03885_ _03893_ VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__nand2_1
X_08938_ _02850_ _00646_ _01536_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__a21o_1
X_08869_ _02781_ _02571_ _00586_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__a21oi_1
X_10900_ _04415_ Qset\[2\]\[11\] VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__nand2_1
X_11880_ _05315_ _05316_ _05703_ _05733_ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__a31o_1
XFILLER_0_67_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10831_ _04042_ _04730_ _04732_ _04734_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_39_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10762_ _04657_ _04659_ _04663_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12501_ _06217_ _06258_ VGND VGND VPWR VPWR _06218_ sky130_fd_sc_hd__nand2_4
X_12432_ _06163_ _06166_ _02125_ VGND VGND VPWR VPWR _00424_ sky130_fd_sc_hd__o21a_1
X_10693_ _04596_ _04597_ VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12363_ _06103_ _06109_ _02125_ VGND VGND VPWR VPWR _00412_ sky130_fd_sc_hd__o21a_1
X_12294_ _06055_ result_reg_set\[3\] VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__nand2_1
X_11314_ _05214_ _05208_ VGND VGND VPWR VPWR _05216_ sky130_fd_sc_hd__nand2_1
X_11245_ _04303_ _05143_ _05144_ _05145_ _05146_ VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__o32a_2
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11176_ _05078_ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__inv_2
X_10127_ _04032_ _03956_ _04033_ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__nand3_1
X_10058_ _03019_ _03876_ VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09910_ _03157_ Qset\[0\]\[8\] VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09841_ _03747_ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06984_ _01102_ _01103_ _00643_ VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__mux2_1
X_09772_ _03678_ _03679_ VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__nand2_1
X_08723_ _02624_ _02146_ VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08654_ _02567_ _02152_ _02560_ _02568_ VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__o211ai_1
X_07605_ _01666_ _00551_ _01282_ _01667_ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__o2bb2a_1
X_08585_ _02470_ _02500_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__nor2_1
X_07536_ _01600_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_105_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09206_ _02529_ _02277_ VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07467_ _01533_ VGND VGND VPWR VPWR _00092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07398_ _01192_ _01463_ _01464_ _01220_ _01470_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__a311o_1
X_06418_ _00552_ VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__buf_2
X_06349_ _00490_ _00484_ VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__nor2_1
X_09137_ _03047_ VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__inv_2
X_09068_ _00622_ _02963_ _02979_ VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08019_ Oset\[1\]\[3\] _01314_ _02019_ VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11030_ _04931_ _04928_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__nand2_1
X_12981_ clknet_leaf_2_clk _00424_ VGND VGND VPWR VPWR CMD_setloop sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11932_ _03122_ _05745_ _03141_ _05749_ _05778_ VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__a221o_2
X_11863_ _05722_ VGND VGND VPWR VPWR _00299_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ _04717_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11794_ _02828_ _02830_ _05673_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10745_ _04507_ _04502_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10676_ _04579_ _04580_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_23_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12415_ _06152_ _06153_ _02116_ VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12346_ im_reg\[9\] net34 _01146_ VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12277_ _06032_ _01075_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11228_ _05128_ _05130_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11159_ _03206_ _03685_ _03697_ _03695_ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__o31a_1
XFILLER_0_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08370_ _02291_ _02294_ VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__nand2_2
XFILLER_0_105_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07321_ _01396_ _01299_ _01208_ _01397_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__a211o_1
XFILLER_0_85_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07252_ Oset\[3\]\[4\] _01332_ _01250_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_07183_ _01264_ VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__buf_2
XFILLER_0_14_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09824_ _03730_ _03731_ _03727_ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__nand3_1
X_06967_ _01086_ _00745_ VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__or2_1
X_09755_ _03662_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__inv_2
X_06898_ net4 _00600_ _00739_ VGND VGND VPWR VPWR _01021_ sky130_fd_sc_hd__a21oi_1
X_09686_ _03591_ VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__inv_2
X_08706_ _02620_ _02577_ VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__nand2_2
XFILLER_0_96_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08637_ _02551_ VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__buf_2
XFILLER_0_68_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08568_ _02470_ Oset\[3\]\[14\] _02374_ _02484_ VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07519_ _01583_ VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08499_ _02415_ _02418_ VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__nand2_2
X_10530_ _03752_ _03755_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10461_ _04151_ _04140_ _04138_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__o21bai_1
X_12200_ result_reg_or\[7\] _05959_ _05992_ _05995_ _05940_ VGND VGND VPWR VPWR _00363_
+ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_20_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10392_ _04297_ _01156_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__nand2_1
X_12131_ _01578_ _04107_ VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12062_ _01209_ _05873_ _05775_ _05880_ VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__a211oi_1
X_11013_ _04915_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12964_ clknet_leaf_6_clk _00407_ VGND VGND VPWR VPWR im_reg\[6\] sky130_fd_sc_hd__dfxtp_4
X_11915_ _05763_ _05743_ VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12895_ clknet_leaf_24_clk _00338_ VGND VGND VPWR VPWR result_reg_Rshift\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_82_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _05706_ _02860_ VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11777_ _05660_ _05661_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10728_ _04610_ _04611_ _04632_ VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__nand3_2
XFILLER_0_70_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10659_ _04537_ _04563_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_93_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12329_ result_reg_set\[15\] _06063_ _06066_ _06084_ VGND VGND VPWR VPWR _00403_
+ sky130_fd_sc_hd__o211a_1
X_07870_ _01093_ _01083_ _01544_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__mux2_1
X_06821_ _00929_ _00725_ _00946_ VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__o21a_1
X_06752_ result_reg_mac\[7\] VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__inv_2
X_09540_ _02653_ _03449_ VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09471_ _03207_ _03211_ _03210_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__a21boi_2
X_06683_ _00541_ _00812_ _00535_ VGND VGND VPWR VPWR _00813_ sky130_fd_sc_hd__a21oi_1
X_08422_ _02329_ _02342_ _02343_ _02344_ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_86_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08353_ _02241_ Oset\[1\]\[5\] _02143_ _02278_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__a211o_1
X_07304_ _01381_ _01238_ _01215_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08284_ _02209_ _02212_ _01551_ VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_34_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07235_ result_reg_Lshift\[4\] result_reg_Rshift\[4\] _01165_ VGND VGND VPWR VPWR
+ _01316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07166_ Oset\[3\]\[0\] _01218_ _01250_ VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__mux2_1
X_07097_ _01181_ VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09807_ Oset\[1\]\[7\] _03033_ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__nand2_1
X_07999_ Oset\[0\]\[10\] _01437_ _02000_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__mux2_1
X_09738_ H\[1\]\[7\] _03341_ _03004_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09669_ _03021_ Oset\[0\]\[6\] VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11700_ Oset\[2\]\[15\] Oset\[3\]\[15\] _03793_ VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__mux2_1
X_12680_ clknet_leaf_1_clk _00130_ VGND VGND VPWR VPWR LC\[4\] sky130_fd_sc_hd__dfxtp_1
X_11631_ _03746_ _05530_ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11562_ _05461_ _05462_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10513_ _02377_ _04415_ _04418_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11493_ _05391_ _05392_ _05393_ VGND VGND VPWR VPWR _05394_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10444_ _04348_ _04349_ VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__nand2_1
X_10375_ _04216_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12114_ _01200_ _04288_ _03846_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__or3_1
X_12045_ _05834_ _05851_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12947_ clknet_leaf_15_clk _00390_ VGND VGND VPWR VPWR result_reg_set\[2\] sky130_fd_sc_hd__dfxtp_1
X_12878_ clknet_leaf_25_clk _00321_ VGND VGND VPWR VPWR result_reg_Lshift\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_160 R2\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11829_ result_reg_mul\[14\] _05677_ _01149_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__o21a_1
XANTENNA_171 _01332_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 _03136_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07020_ _01124_ VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08971_ _02873_ _01154_ _02882_ VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__nand3_1
X_07922_ Oset\[2\]\[14\] _01508_ _01941_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__mux2_1
X_07853_ net6 _01746_ VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__nor2_1
X_06804_ result_reg_set\[9\] VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__inv_2
X_07784_ _01835_ _01838_ _01612_ VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_67_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06735_ _00553_ result_reg_or\[6\] VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__or2b_1
X_09523_ Qset\[3\]\[5\] _03024_ _02837_ VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__a21oi_1
X_06666_ result_reg_sub\[4\] _00740_ _00796_ VGND VGND VPWR VPWR _00797_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_66_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09454_ _03361_ VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__inv_2
X_09385_ _03295_ VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08405_ _02250_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__clkbuf_4
X_06597_ _00611_ VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__buf_4
X_08336_ _02260_ H\[1\]\[4\] _02262_ VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__o21ai_1
X_08267_ _02127_ Qset\[3\]\[2\] VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__nand2_1
X_07218_ result_reg_and\[3\] _01299_ VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08198_ _02128_ VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__buf_6
X_07149_ shift.left CMD_logic_shift_right _00624_ _01233_ VGND VGND VPWR VPWR _01234_
+ sky130_fd_sc_hd__or4_1
XFILLER_0_61_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10160_ _02565_ H\[0\]\[14\] VGND VGND VPWR VPWR _04067_ sky130_fd_sc_hd__nor2_1
X_10091_ _03996_ _03964_ _03968_ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12801_ clknet_leaf_10_clk _00244_ VGND VGND VPWR VPWR result_reg_add\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10993_ _04895_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__inv_4
X_12732_ clknet_leaf_37_clk _00175_ VGND VGND VPWR VPWR H\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_12663_ clknet_3_0__leaf_clk _00113_ VGND VGND VPWR VPWR Oset\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_11614_ _04302_ H\[2\]\[15\] _05513_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__a21o_1
X_12594_ clknet_leaf_48_clk _00044_ VGND VGND VPWR VPWR Qset\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11545_ _05439_ _05445_ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__or2_1
X_11476_ _05253_ _05248_ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__nand2_1
X_10427_ _04328_ _04332_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_90_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10358_ _04210_ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10289_ _03897_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_29_Left_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12028_ _01148_ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06520_ _00654_ VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06451_ shift.H VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__buf_6
XFILLER_0_8_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06382_ im_reg\[8\] _00486_ VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09170_ _02528_ _02292_ VGND VGND VPWR VPWR _03081_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08121_ H\[0\]\[2\] _01676_ _02075_ VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08052_ _01676_ H\[2\]\[2\] _02038_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__mux2_1
X_07003_ _00878_ Qset\[1\]\[6\] _01109_ VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_47_Left_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08954_ _02864_ _02525_ _02865_ VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__nand3_1
X_07905_ _01948_ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__clkbuf_1
X_08885_ _02561_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__buf_6
XFILLER_0_98_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07836_ _01586_ result_reg_sub\[13\] VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__nand2_1
X_07767_ result_reg_mul\[10\] _01679_ _01656_ VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06718_ _00811_ _00695_ _00836_ _00847_ _00644_ VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_56_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09506_ _03373_ _03377_ _03274_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__nand3_1
XFILLER_0_39_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07698_ _01756_ result_reg_mac\[6\] _01570_ VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__mux2_1
X_06649_ result_reg_Rshift\[3\] _00753_ _00780_ VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__o21ai_1
X_09437_ _03346_ _02572_ _00587_ VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__a21oi_1
X_09368_ _03277_ _03278_ VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08319_ _02244_ _02147_ _02245_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__nand3_1
X_09299_ _03200_ _03203_ VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_82 _01712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 _01485_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11330_ _05079_ _04309_ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__nor2_1
XANTENNA_60 _01368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 _01801_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11261_ _05159_ _05160_ _05161_ _05162_ _00621_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_76_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13000_ clknet_leaf_39_clk _00443_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dfxtp_1
X_11192_ _04308_ _04651_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__nand2_1
X_10212_ _04116_ _04100_ _04101_ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_100_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10143_ _04049_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__inv_2
X_10074_ _03980_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_74_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10976_ _04878_ _03274_ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12715_ clknet_leaf_44_clk _00158_ VGND VGND VPWR VPWR Oset\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12646_ clknet_leaf_49_clk _00096_ VGND VGND VPWR VPWR H\[3\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_562 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12577_ clknet_leaf_48_clk _00027_ VGND VGND VPWR VPWR Qset\[0\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11528_ _05427_ _05413_ VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11459_ _05243_ _05232_ _05242_ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08670_ _02579_ VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__buf_6
X_07621_ _01306_ _01682_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_49_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07552_ _00670_ _01593_ VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__nor2_1
X_06503_ _00623_ _00557_ VGND VGND VPWR VPWR _00638_ sky130_fd_sc_hd__nor2_1
X_07483_ _01547_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__inv_2
X_06434_ _00568_ VGND VGND VPWR VPWR _00569_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09222_ _03132_ VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06365_ _00503_ _00475_ _00504_ next_PC\[5\] _00478_ VGND VGND VPWR VPWR _00019_
+ sky130_fd_sc_hd__a32o_1
X_09153_ _03063_ _02552_ VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__nand2_1
X_08104_ _02068_ VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__clkbuf_1
X_06296_ _06261_ current_state\[1\] VGND VGND VPWR VPWR _06262_ sky130_fd_sc_hd__or2b_1
X_09084_ _02582_ Qset\[0\]\[4\] VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__nand2_1
X_08035_ Oset\[1\]\[11\] _01455_ _02018_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09986_ _03892_ VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__inv_2
X_08937_ _02837_ _02847_ _02849_ VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__o21ai_1
X_08868_ _02778_ _02780_ VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__nand2_2
X_07819_ result_reg_or\[12\] _01595_ _01593_ VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__o21ai_1
X_08799_ _02712_ VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10830_ _04729_ Oset\[3\]\[11\] _04045_ _04733_ VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10761_ _04660_ _04664_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12500_ _06216_ _06266_ _06263_ VGND VGND VPWR VPWR _06217_ sky130_fd_sc_hd__and3_1
X_10692_ _04595_ _04571_ _04572_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_94_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12431_ _06165_ _06160_ VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__nor2_1
X_12362_ _06105_ _06106_ _06102_ _06108_ VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_10_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12293_ _06058_ R2\[1\] VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__nand2_1
X_11313_ _05208_ _05214_ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11244_ Qset\[1\]\[13\] _04302_ _04303_ VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__o21ai_1
X_11175_ _03897_ _03206_ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__nor2_1
X_10126_ _03922_ _03944_ VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__and2_1
X_10057_ _03930_ _03963_ VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10959_ _03798_ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12629_ clknet_leaf_45_clk _00079_ VGND VGND VPWR VPWR Oset\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ _03744_ _03746_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06983_ result_reg_Lshift\[15\] VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__inv_2
X_09771_ _03667_ _03668_ _03671_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__nand3_1
X_08722_ Oset\[3\]\[0\] _02624_ _02626_ _02636_ VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08653_ H\[3\]\[0\] _02567_ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__nand2_1
X_07604_ _01588_ VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__clkbuf_4
X_08584_ Qset\[2\]\[15\] VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__inv_2
X_07535_ _00921_ _01556_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__nor2_4
XFILLER_0_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07466_ _01531_ _01532_ VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06417_ _00551_ _00526_ VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__nand2_2
XFILLER_0_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09205_ _03051_ _03115_ VGND VGND VPWR VPWR _03116_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07397_ net4 _01187_ _01254_ _01469_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__o211a_1
X_06348_ next_PC\[3\] VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09136_ _00583_ _02551_ VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09067_ _01536_ _02965_ _02967_ _00549_ _02978_ VGND VGND VPWR VPWR _02979_ sky130_fd_sc_hd__a311o_1
X_08018_ _02022_ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_73_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09969_ _03875_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__buf_4
X_12980_ clknet_leaf_3_clk _00423_ VGND VGND VPWR VPWR CMD_loopjump sky130_fd_sc_hd__dfxtp_1
X_11931_ _00591_ _05777_ VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__nor2_1
X_11862_ _00880_ _05707_ _05710_ _05721_ VGND VGND VPWR VPWR _05722_ sky130_fd_sc_hd__a211o_1
XFILLER_0_86_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10813_ _04714_ _04716_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11793_ result_reg_mul\[1\] _05670_ _05672_ _05674_ VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_476 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10744_ _03701_ _03703_ VGND VGND VPWR VPWR _04648_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10675_ _04074_ _03020_ _04096_ _02963_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_23_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12414_ _06126_ CMD_load VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__nand2_1
X_12345_ _06094_ VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12276_ _06039_ _05828_ _06044_ _06049_ VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11227_ _05129_ _05120_ VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__nand2_1
X_11158_ _03701_ _03699_ VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__nand2_1
X_10109_ _04014_ _04015_ VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__nand2_1
X_11089_ _04691_ _04899_ _04991_ VGND VGND VPWR VPWR _04992_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_59_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07320_ _00559_ result_reg_and\[8\] _01243_ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07251_ _01161_ _01317_ _01331_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__a21bo_4
XTAP_TAPCELL_ROW_98_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07182_ _01265_ VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09823_ _03705_ _00831_ _03706_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__nand3_1
XFILLER_0_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06966_ result_reg_mul\[15\] VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__inv_2
X_09754_ _03660_ _03508_ _03661_ VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__a21oi_1
X_06897_ result_reg_set\[12\] _00615_ _00696_ _01019_ VGND VGND VPWR VPWR _01020_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_55_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09685_ _03571_ _02092_ _03572_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__nand3_1
X_08705_ _02619_ VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__buf_6
X_08636_ _02539_ VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__inv_2
X_08567_ _02470_ _02483_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07518_ _01578_ _00533_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__nor2_2
XFILLER_0_49_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08498_ _02364_ Oset\[1\]\[11\] _02329_ _02417_ VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__a211o_1
X_07449_ _01086_ _01518_ _01177_ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10460_ _04040_ _04365_ _04028_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__nand3_1
XFILLER_0_44_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09119_ H\[1\]\[4\] _03025_ _02840_ VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10391_ _03770_ _04288_ _04296_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12130_ _01243_ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__clkbuf_4
X_12061_ _05875_ _05877_ _05878_ _05879_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11012_ _04913_ _04914_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__nand2_1
X_12963_ clknet_3_1__leaf_clk _00406_ VGND VGND VPWR VPWR R1\[1\] sky130_fd_sc_hd__dfxtp_4
X_11914_ _05759_ _05762_ _05755_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ clknet_leaf_24_clk _00337_ VGND VGND VPWR VPWR result_reg_Rshift\[13\] sky130_fd_sc_hd__dfxtp_1
X_11845_ _00635_ VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__buf_4
XFILLER_0_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11776_ _05628_ _01067_ _02650_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10727_ _04630_ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__inv_2
X_10658_ _04561_ _04562_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10589_ _04493_ _02403_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__nand2_8
XTAP_TAPCELL_ROW_93_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12328_ im_reg\[7\] _05745_ R2\[1\] _05744_ _06054_ VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__a221o_1
X_12259_ _06039_ _05779_ _06013_ _06040_ VGND VGND VPWR VPWR _00377_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_10_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06820_ _00938_ _00619_ _00629_ _00945_ VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__a211o_1
XFILLER_0_92_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06751_ _00879_ VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__clkbuf_1
X_06682_ result_reg_add\[5\] VGND VGND VPWR VPWR _00812_ sky130_fd_sc_hd__inv_2
X_09470_ _03228_ _03216_ _03214_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__o21bai_1
X_08421_ Oset\[1\]\[8\] _02260_ _02254_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08352_ _02141_ _02277_ VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__nor2_1
X_07303_ _01377_ _01380_ _00890_ _01271_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_58_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08283_ _02151_ _02210_ _00003_ _02211_ VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_34_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07234_ _01315_ VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07165_ _01249_ VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__buf_4
X_07096_ _01179_ _01180_ VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__nand2_4
XFILLER_0_41_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09806_ _03021_ Oset\[0\]\[7\] VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__nand2_1
X_07998_ _02011_ VGND VGND VPWR VPWR _00145_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06949_ _01066_ _01069_ _00608_ VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__mux2_1
X_09737_ _03498_ H\[0\]\[7\] VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__nor2_1
X_09668_ H\[1\]\[6\] _03025_ _02840_ _03576_ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_25_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ _02533_ VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__buf_6
X_09599_ _03507_ _03258_ VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__nor2_1
X_11630_ _05528_ _05529_ VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11561_ _05460_ _05456_ _05457_ VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_92_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10512_ _04415_ H\[0\]\[9\] _03798_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__a21oi_1
X_11492_ _05268_ _05257_ _05267_ VGND VGND VPWR VPWR _05393_ sky130_fd_sc_hd__a21o_1
X_10443_ _03506_ _03868_ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_79_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10374_ _04277_ _04279_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12113_ _05922_ _05803_ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__nand2_1
X_12044_ _05866_ VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12946_ clknet_leaf_15_clk _00389_ VGND VGND VPWR VPWR result_reg_set\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12877_ clknet_leaf_25_clk _00320_ VGND VGND VPWR VPWR result_reg_Lshift\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_161 R3\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_150 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_172 _01362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_183 _05634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11828_ _05697_ VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__inv_2
X_11759_ _05627_ _04444_ VGND VGND VPWR VPWR _05649_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_579 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08970_ _02881_ _02551_ VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__nand2_1
X_07921_ _01956_ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__clkbuf_1
X_07852_ _01066_ _01682_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__or2_1
Xinput1 data_in[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
X_06803_ result_reg_mac\[9\] VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__inv_2
X_07783_ result_reg_not\[10\] _01633_ _01837_ VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_67_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09522_ Qset\[1\]\[5\] _03024_ VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_48_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_39_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06734_ _00859_ _00743_ _00861_ _00862_ VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__a31o_1
X_06665_ _00540_ _00789_ _00534_ VGND VGND VPWR VPWR _00796_ sky130_fd_sc_hd__a21oi_1
X_09453_ _03270_ _03265_ _03264_ VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__a21oi_1
X_09384_ _00789_ _02654_ _02753_ _03294_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__a211o_1
X_08404_ _02261_ VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__buf_4
X_06596_ result_reg_add\[2\] VGND VGND VPWR VPWR _00729_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08335_ _02261_ H\[0\]\[4\] _02254_ VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08266_ _02128_ Qset\[2\]\[2\] VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__nand2_1
X_07217_ _01207_ VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__clkbuf_4
X_08197_ _02127_ VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__inv_6
X_07148_ CMD_not _00545_ CMD_and _01232_ VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07079_ _01163_ _00641_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__nand2_4
X_10090_ _03964_ _03968_ _03996_ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_39_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
X_12800_ clknet_leaf_39_clk _00243_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10992_ _04893_ _04894_ VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_2_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ clknet_leaf_41_clk _00174_ VGND VGND VPWR VPWR H\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12662_ clknet_leaf_45_clk _00112_ VGND VGND VPWR VPWR Oset\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_11613_ _05335_ H\[3\]\[15\] _04303_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12593_ clknet_leaf_48_clk _00043_ VGND VGND VPWR VPWR Qset\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11544_ _05443_ _05444_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__and2_1
X_11475_ _05374_ _05375_ VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__nand2_1
X_10426_ _04331_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10357_ _04219_ _04214_ _04213_ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__a21boi_1
X_10288_ _04193_ _04194_ _03751_ VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__a21o_1
X_12027_ result_reg_Rshift\[5\] _05848_ _05808_ _05856_ VGND VGND VPWR VPWR _00329_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12929_ clknet_leaf_19_clk _00372_ VGND VGND VPWR VPWR result_reg_not\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06450_ _00584_ VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__buf_4
X_06381_ _00516_ _00517_ _00486_ VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_71_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08120_ _02077_ VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08051_ _02040_ VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__clkbuf_1
X_07002_ _01115_ VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08953_ _02544_ Qset\[3\]\[3\] VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07904_ Oset\[2\]\[5\] _01349_ _01942_ VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__mux2_1
X_08884_ _02794_ _02796_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__nand2_1
X_07835_ _01581_ result_reg_add\[13\] VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__nand2_1
X_07766_ _00958_ _00959_ _01545_ VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__mux2_1
X_06717_ _00650_ _00846_ VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09505_ _03413_ _02092_ _03414_ VGND VGND VPWR VPWR _03415_ sky130_fd_sc_hd__nand3_1
X_07697_ _01594_ _01748_ _01755_ VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__o21ai_1
X_09436_ _03342_ _03343_ _03344_ _03345_ VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__a22oi_4
X_06648_ _00754_ _00779_ VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__nand2_1
X_06579_ _00557_ _00631_ _00634_ _00712_ VGND VGND VPWR VPWR _00713_ sky130_fd_sc_hd__or4_1
X_09367_ _03206_ _00549_ VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__nand2_1
XANTENNA_50 _01205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08318_ _02141_ Qset\[1\]\[4\] VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__nand2_1
X_09298_ _03202_ _03204_ _03208_ VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__nand3_1
XFILLER_0_105_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_83 _01714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 _01380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _01488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08249_ Oset\[2\]\[1\] VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_94 _01801_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11260_ Qset\[1\]\[13\] _04857_ VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10211_ _02949_ _04110_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__nor2_1
X_11191_ _04494_ _04460_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10142_ _03758_ _04048_ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__nor2_2
XFILLER_0_30_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10073_ _03938_ _03935_ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10975_ _04825_ _04877_ _04824_ VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__nand3_1
X_12714_ clknet_leaf_45_clk _00157_ VGND VGND VPWR VPWR Oset\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12645_ clknet_leaf_53_clk _00095_ VGND VGND VPWR VPWR H\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12576_ clknet_leaf_45_clk _00026_ VGND VGND VPWR VPWR Qset\[0\]\[2\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_13_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11527_ _05413_ _05427_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11458_ _05288_ _05280_ VGND VGND VPWR VPWR _05359_ sky130_fd_sc_hd__nand2_1
X_11389_ _04176_ _05290_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__xor2_1
X_10409_ _04314_ _04263_ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07620_ _01560_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_49_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07551_ R1\[1\] _01541_ _01606_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__o21a_1
X_06502_ CMD_logic_shift_right VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__inv_2
X_07482_ _01542_ _00533_ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06433_ _00567_ _00538_ VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__nor2_2
XFILLER_0_63_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09221_ _02556_ _03131_ VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09152_ _03060_ _03062_ VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__nand2_2
X_06364_ R1\[1\] _00486_ VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08103_ _01839_ H\[1\]\[10\] _02056_ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06295_ _06258_ _06259_ VGND VGND VPWR VPWR _06261_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_2_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09083_ _02990_ _02991_ _02993_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__nand3_1
X_08034_ _02030_ VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09985_ _03886_ _03891_ _03888_ VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__o21ai_1
X_08936_ Qset\[0\]\[2\] _02632_ _02848_ VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__a21o_1
X_08867_ _02586_ H\[1\]\[2\] _02584_ _02779_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__a211o_1
X_07818_ _01691_ result_reg_and\[12\] VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__nand2_1
X_08798_ _00580_ _00669_ _02539_ VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__o21ai_1
X_07749_ _01804_ result_reg_mul\[9\] _01583_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10760_ _04663_ VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__inv_2
X_10691_ _04573_ _04595_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__nand2_1
X_09419_ _03328_ _00581_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__nand2_1
X_12430_ _06115_ _06164_ VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12361_ _06107_ _06100_ _06253_ _06098_ VGND VGND VPWR VPWR _06108_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_10_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12292_ _06059_ _06060_ _02116_ VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__a21oi_1
X_11312_ _05209_ _05213_ VGND VGND VPWR VPWR _05214_ sky130_fd_sc_hd__xnor2_1
X_11243_ _04832_ Qset\[0\]\[13\] VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11174_ _03206_ _05063_ _05076_ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__or3_1
XFILLER_0_38_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10125_ _03984_ _04008_ VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__nor2_1
X_10056_ _03019_ _03868_ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_46_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10958_ H\[2\]\[12\] _04856_ _04860_ VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10889_ _04744_ _02096_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__nand2_1
X_12628_ clknet_leaf_43_clk _00078_ VGND VGND VPWR VPWR Oset\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12559_ _06250_ VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06982_ result_reg_Rshift\[15\] VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__inv_2
X_09770_ _03669_ _03673_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__nand2_1
X_08721_ _02624_ _02142_ VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__nor2_1
X_08652_ _02529_ VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__buf_6
X_07603_ _01571_ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08583_ _02499_ VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__clkbuf_1
X_07534_ result_reg_mac\[0\] _01541_ _01598_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_105_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07465_ _00472_ VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_93_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06416_ _00530_ _00545_ _00528_ _00550_ VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__and4_2
X_09204_ _02784_ VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07396_ _01468_ _01187_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06347_ R2\[1\] _06285_ VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__or2_1
X_09135_ _00624_ _03020_ _03045_ VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_102_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09066_ _02972_ _02977_ _01536_ VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_558 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08017_ Oset\[1\]\[2\] _01295_ _02019_ VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09968_ _03874_ _01552_ _02572_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__and3_1
X_08919_ _02821_ _00549_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__nand2_1
X_11930_ _03128_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__inv_2
X_09899_ Qset\[2\]\[8\] _03025_ VGND VGND VPWR VPWR _03806_ sky130_fd_sc_hd__or2_1
X_11861_ _05706_ _03740_ VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11792_ _02737_ _02740_ _05673_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_43_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _04709_ _04710_ _04715_ VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__nand3_1
XFILLER_0_67_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10743_ _04514_ _04511_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10674_ _04369_ _04578_ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_23_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12413_ _06266_ _06148_ _06151_ VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__or3b_1
XFILLER_0_35_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12344_ _06093_ _01532_ VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12275_ _06032_ _01049_ VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11226_ _05127_ _04878_ _03274_ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__nand3_1
X_11157_ _04709_ _04702_ VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__nand2_1
X_10108_ _04013_ _03989_ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__nand2_1
X_11088_ _04989_ _04990_ VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_59_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10039_ _03911_ _03945_ VGND VGND VPWR VPWR _03946_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07250_ _01322_ _01215_ _01329_ _01159_ _01330_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_98_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07181_ _01204_ VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09822_ _03707_ _02092_ VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__nand2_1
X_09753_ _03473_ _03471_ VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__nor2_1
X_06965_ result_reg_sub\[15\] _00541_ _01084_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__o21ai_2
X_08704_ _02618_ _02158_ VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__nand2_4
X_06896_ _01018_ _00615_ VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__nand2_1
X_09684_ _03566_ _00536_ _03567_ VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__nand3_1
XFILLER_0_96_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08635_ _02547_ _02549_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__nand2_2
XFILLER_0_96_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08566_ Oset\[2\]\[14\] VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__inv_2
X_07517_ _01581_ result_reg_add\[0\] VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08497_ _02356_ _02416_ VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__nor2_1
X_07448_ _01093_ _01083_ _01174_ VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07379_ _01192_ _01445_ _01446_ _01220_ _01452_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_20_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09118_ H\[2\]\[4\] _03023_ _03028_ VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__a21o_1
X_10390_ _04289_ _04295_ _03770_ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__nand3_1
X_09049_ _02959_ Add.sub VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__nand2_1
X_12060_ _00525_ _02538_ _02595_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__or3_1
X_11011_ _04912_ _04898_ VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__nand2_1
X_12962_ clknet_leaf_52_clk _00405_ VGND VGND VPWR VPWR R2\[1\] sky130_fd_sc_hd__dfxtp_4
X_12893_ clknet_leaf_24_clk _00336_ VGND VGND VPWR VPWR result_reg_Rshift\[12\] sky130_fd_sc_hd__dfxtp_1
X_11913_ _05744_ _05760_ _05761_ VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_56_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _05709_ VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11775_ _05485_ _05486_ _05655_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__nand3_1
X_10726_ _04612_ _04630_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10657_ _04560_ _04538_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10588_ _04492_ _01553_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_93_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12327_ result_reg_set\[14\] _06063_ _06066_ _06083_ VGND VGND VPWR VPWR _00402_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12258_ _06033_ _00849_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__nand2_1
X_11209_ _05111_ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__inv_2
X_12189_ _03091_ _03482_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__nand2_1
X_06750_ _00878_ Qset\[0\]\[6\] _00687_ VGND VGND VPWR VPWR _00879_ sky130_fd_sc_hd__mux2_1
X_06681_ result_reg_mac\[5\] VGND VGND VPWR VPWR _00811_ sky130_fd_sc_hd__inv_2
X_08420_ _02319_ Oset\[0\]\[8\] VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08351_ Oset\[0\]\[5\] VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__inv_2
X_07302_ result_reg_mul\[7\] _01263_ _01245_ _01379_ VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08282_ H\[1\]\[2\] _02129_ VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__nor2_1
X_07233_ Oset\[3\]\[3\] _01314_ _01250_ VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07164_ _01225_ _01248_ VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__nor2_4
X_07095_ _00579_ _00653_ VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07997_ Oset\[0\]\[9\] _01420_ _02001_ VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__mux2_1
X_09805_ H\[0\]\[7\] _03022_ _03712_ VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__a21o_1
X_06948_ _01060_ _01068_ _00613_ VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__mux2_1
X_09736_ H\[2\]\[7\] H\[3\]\[7\] _02611_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__mux2_1
X_09667_ _03025_ _02303_ VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__nor2_1
X_06879_ _00999_ _00655_ _00657_ _01002_ _00666_ VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__a221o_1
X_08618_ _00007_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _03506_ VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_81_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ H\[2\]\[13\] H\[3\]\[13\] _02459_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11560_ _05458_ _05460_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10511_ H\[2\]\[9\] _04415_ _04416_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11491_ _05390_ _05380_ VGND VGND VPWR VPWR _05392_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10442_ _03652_ _03876_ VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_79_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10373_ _04272_ _04275_ _04278_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__nand3_1
X_12112_ _01578_ _04305_ VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12043_ _05829_ _05851_ _05775_ _05865_ VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_5_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12945_ clknet_leaf_14_clk _00388_ VGND VGND VPWR VPWR result_reg_set\[0\] sky130_fd_sc_hd__dfxtp_1
X_12876_ clknet_leaf_24_clk _00319_ VGND VGND VPWR VPWR result_reg_Lshift\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_140 _06218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_151 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_173 _01415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_184 _05634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11827_ _05229_ _05298_ _05677_ _05696_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_162 R3\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11758_ _05648_ VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10709_ H\[2\]\[10\] _04414_ _04613_ VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11689_ _05558_ _05588_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__xor2_1
XFILLER_0_70_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07920_ Oset\[2\]\[13\] _01490_ _01941_ VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__mux2_1
X_07851_ _01900_ _01653_ _01901_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__a21o_1
Xinput2 data_in[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dlymetal6s2s_1
X_07782_ result_reg_Rshift\[10\] _01672_ _01607_ _01836_ VGND VGND VPWR VPWR _01837_
+ sky130_fd_sc_hd__o211a_1
X_06802_ _00928_ VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__clkbuf_1
X_06733_ result_reg_and\[6\] _00743_ _00553_ VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_67_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09521_ _02632_ Qset\[0\]\[5\] VGND VGND VPWR VPWR _03431_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_39_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06664_ result_reg_or\[4\] VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09452_ _03300_ _03361_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__nand2_1
X_09383_ _02653_ _03293_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__nor2_1
X_06595_ result_reg_sub\[2\] VGND VGND VPWR VPWR _00728_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08403_ _02260_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__clkbuf_4
X_08334_ _02141_ VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__buf_4
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08265_ _02194_ VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__clkbuf_1
X_07216_ result_reg_not\[3\] _01297_ _01168_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08196_ _00002_ VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__buf_6
X_07147_ _01157_ CMD_set VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07078_ _01162_ _00531_ VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__nor2_2
X_10991_ _04108_ _03745_ VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09719_ _03626_ _03610_ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12730_ clknet_leaf_44_clk _00173_ VGND VGND VPWR VPWR H\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_12661_ clknet_leaf_53_clk _00111_ VGND VGND VPWR VPWR Oset\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11612_ _05511_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__inv_2
X_12592_ clknet_leaf_46_clk _00042_ VGND VGND VPWR VPWR Qset\[1\]\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_92_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11543_ _05441_ _05440_ VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__nand2_1
X_11474_ _05373_ _05360_ VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__nand2_1
X_10425_ _03950_ _04330_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10356_ _04234_ _04261_ VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10287_ _04192_ _04159_ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__nand2_1
X_12026_ _05786_ _05851_ VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12928_ clknet_leaf_16_clk _00371_ VGND VGND VPWR VPWR result_reg_or\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_36_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ clknet_leaf_18_clk _00302_ VGND VGND VPWR VPWR result_reg_mac\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06380_ _00511_ _00515_ VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08050_ _01650_ H\[2\]\[1\] _02038_ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07001_ _00854_ Qset\[1\]\[5\] _01109_ VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08952_ _02787_ Qset\[2\]\[3\] VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__nand2_1
X_08883_ _02795_ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__inv_2
X_07903_ _01947_ VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__clkbuf_1
X_07834_ _01883_ _01658_ _01884_ _01885_ VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__a31o_1
X_07765_ _01820_ VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__clkbuf_1
X_07696_ _01752_ _01572_ _01753_ _01568_ _01754_ VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__a311o_1
X_06716_ net12 _00735_ _00839_ _00845_ VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__o211a_1
X_09504_ _03145_ _00556_ VGND VGND VPWR VPWR _03414_ sky130_fd_sc_hd__nand2_1
X_06647_ result_reg_Lshift\[3\] VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__inv_2
X_09435_ _02991_ VGND VGND VPWR VPWR _03345_ sky130_fd_sc_hd__buf_4
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06578_ shift.left CMD_logic_shift_right _00710_ _00711_ VGND VGND VPWR VPWR _00712_
+ sky130_fd_sc_hd__or4_1
X_09366_ _03234_ _03276_ _00622_ VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__nand3_1
XANTENNA_40 _01044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08317_ _02230_ Qset\[0\]\[4\] VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__nand2_1
X_09297_ _03207_ VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_84 _01727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 _01496_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 _01396_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 _01270_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08248_ _02174_ _02177_ VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__nand2_2
XFILLER_0_34_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_95 _01806_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08179_ im_reg\[8\] _02100_ _02105_ _02113_ VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__o211a_1
X_10210_ _04102_ _04116_ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_76_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11190_ _04494_ _04651_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__nand2_1
X_10141_ _00588_ _04047_ VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_7_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10072_ _03976_ _03978_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10974_ _04816_ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_43_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12713_ clknet_leaf_44_clk _00156_ VGND VGND VPWR VPWR Oset\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12644_ clknet_leaf_49_clk _00094_ VGND VGND VPWR VPWR H\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12575_ clknet_leaf_46_clk _00025_ VGND VGND VPWR VPWR Qset\[0\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11526_ _05426_ VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11457_ _05296_ _05293_ VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11388_ _04177_ _04172_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__or2b_1
X_10408_ _04311_ _04312_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10339_ _04245_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12009_ _05843_ VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07550_ _01599_ _01606_ _01614_ VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06501_ _00635_ _00605_ VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__nor2_2
X_07481_ _00610_ _00542_ _01545_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09220_ _00583_ R1\[1\] VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__nand2_1
X_06432_ _00533_ _00566_ VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09151_ _02874_ Oset\[1\]\[7\] _02727_ _03061_ VGND VGND VPWR VPWR _03062_ sky130_fd_sc_hd__a211o_1
X_06363_ _00501_ _00502_ _00486_ VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_29_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08102_ _02067_ VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09082_ _02992_ Qset\[3\]\[4\] VGND VGND VPWR VPWR _02993_ sky130_fd_sc_hd__nand2_1
X_06294_ net35 _06258_ _06260_ VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08033_ Oset\[1\]\[10\] _01437_ _02018_ VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__mux2_1
X_09984_ _03888_ _03890_ VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__nand2_1
X_08935_ Qset\[1\]\[2\] _02625_ _00001_ VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__a21o_1
X_08866_ _02592_ _02210_ VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07817_ _01867_ _01585_ _01868_ _01869_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__a31o_1
X_08797_ _02707_ _02710_ VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_103_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07748_ result_reg_add\[9\] result_reg_sub\[9\] _01579_ VGND VGND VPWR VPWR _01804_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07679_ result_reg_not\[5\] _01633_ _01738_ VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10690_ _04593_ _04594_ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__nand2_1
X_09418_ _03322_ _03324_ _03327_ VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__o21ai_2
X_09349_ _03256_ _03259_ VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12360_ net22 net21 VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11311_ _05211_ _05212_ VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_10_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12291_ _06055_ result_reg_set\[2\] VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11242_ Qset\[3\]\[13\] _04302_ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__nor2_1
X_11173_ _05074_ _05075_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__nand2_1
X_10124_ _04010_ _04007_ _04030_ VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_89_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10055_ _03858_ _03050_ _03421_ VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_46_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10957_ H\[3\]\[12\] _04858_ _04859_ VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__a21o_1
X_10888_ _04722_ _04791_ _00820_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__nand3_1
X_12627_ clknet_3_0__leaf_clk _00077_ VGND VGND VPWR VPWR Oset\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12558_ _01106_ Qset\[3\]\[15\] _06233_ VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12489_ _06210_ VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__clkbuf_1
X_11509_ _05407_ _05296_ _05293_ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__nand3_1
XFILLER_0_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06981_ result_reg_not\[15\] VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__inv_2
X_08720_ _02626_ _02631_ _02634_ VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__o21a_1
X_08651_ _02565_ _02155_ VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__nor2_1
X_07602_ _01661_ _01585_ _01662_ _01664_ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__a31o_1
X_08582_ _02498_ net53 _02169_ VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__mux2_1
X_07533_ _01565_ _01569_ _01570_ _01597_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__a211o_1
XFILLER_0_44_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07464_ _00498_ net29 current_state\[2\] VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06415_ _00546_ _00547_ _00549_ VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__and3_2
XFILLER_0_63_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09203_ _03109_ _03113_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__nand2_1
X_07395_ _01465_ _01467_ _01182_ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09134_ _01537_ _03029_ _03031_ _00556_ _03044_ VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__a311o_2
X_06346_ _00487_ _00475_ _00488_ next_PC\[2\] _00478_ VGND VGND VPWR VPWR _00016_
+ sky130_fd_sc_hd__a32o_1
X_09065_ _02973_ _02974_ _02975_ _02976_ _00646_ VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08016_ _02021_ VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_73_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09967_ _03870_ _03871_ _02800_ _03872_ _03873_ VGND VGND VPWR VPWR _03874_ sky130_fd_sc_hd__a32o_2
X_08918_ _02828_ _02830_ _00622_ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__nand3_1
X_09898_ Qset\[0\]\[8\] Qset\[1\]\[8\] _03791_ VGND VGND VPWR VPWR _03805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08849_ _02201_ _02161_ VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__nand2_1
X_11860_ _05720_ VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_84_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11791_ _05669_ VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_43_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _04713_ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10742_ _04526_ _04645_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10673_ _04096_ _03020_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__nand2_1
X_12412_ _06150_ net25 VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_51_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12343_ im_reg\[8\] net33 _01146_ VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12274_ _06039_ _05821_ _06044_ _06048_ VGND VGND VPWR VPWR _00384_ sky130_fd_sc_hd__o211a_1
X_11225_ _04880_ _05121_ _05127_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__nand3_1
XFILLER_0_31_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11156_ _05058_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__inv_2
X_11087_ _04988_ _04979_ VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__nand2_1
X_10107_ _03989_ _04013_ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__or2_1
X_10038_ _03910_ VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_59_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11989_ _05827_ VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07180_ _01202_ VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09821_ _03708_ _03709_ _03728_ VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__nand3_1
X_09752_ _03471_ _03473_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__nand2_1
X_06964_ _00740_ _01083_ _00535_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__a21oi_1
X_08703_ _02617_ _01551_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__nand2_1
X_06895_ _01010_ _01017_ _00732_ VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__mux2_1
X_09683_ _03568_ _03573_ _03591_ VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__nand3_1
X_08634_ _02545_ _02146_ _02535_ _02548_ VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_89_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08565_ _02478_ _02481_ VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__nand2_2
X_07516_ _01580_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__clkbuf_4
X_08496_ Oset\[0\]\[11\] VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07447_ result_reg_or\[15\] _01199_ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__or2_1
X_07378_ net3 _01187_ _01254_ _01451_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__o211a_1
X_06329_ _00473_ VGND VGND VPWR VPWR _00474_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09117_ H\[3\]\[4\] _03025_ _03027_ VGND VGND VPWR VPWR _03028_ sky130_fd_sc_hd__a21o_1
X_09048_ Add.sub _02959_ VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11010_ _04898_ _04912_ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12961_ clknet_leaf_54_clk _00404_ VGND VGND VPWR VPWR R3\[1\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_99_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12892_ clknet_leaf_24_clk _00335_ VGND VGND VPWR VPWR result_reg_Rshift\[11\] sky130_fd_sc_hd__dfxtp_1
X_11912_ _01158_ _02881_ _02891_ _05749_ VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_56_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _00694_ _05707_ _05634_ _05708_ VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11774_ _05659_ VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10725_ _00624_ _04494_ _04629_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_82_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10656_ _04538_ _04560_ VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10587_ _04485_ _03758_ _04486_ _04491_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12326_ R2\[0\] _05744_ im_reg\[6\] _05745_ _06054_ VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__a221o_1
X_12257_ _06031_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__buf_2
XFILLER_0_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12188_ result_reg_or\[5\] _05959_ _05983_ _05985_ _05940_ VGND VGND VPWR VPWR _00361_
+ sky130_fd_sc_hd__o221a_1
X_11208_ _05059_ _05110_ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__xor2_1
XFILLER_0_76_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11139_ _05028_ _05041_ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06680_ _00810_ VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__clkbuf_1
X_08350_ _02241_ Oset\[3\]\[5\] _02147_ _02275_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_102_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07301_ result_reg_add\[7\] _01264_ _01266_ _01378_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08281_ H\[0\]\[2\] VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__inv_2
X_07232_ _01161_ _01298_ _01312_ _01313_ VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__a22o_4
XFILLER_0_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07163_ _01242_ _01247_ VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__or2b_2
XFILLER_0_26_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07094_ _00471_ _00558_ _01157_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09804_ H\[1\]\[7\] _03025_ _02840_ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__a21o_1
X_07996_ _02010_ VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__clkbuf_1
X_06947_ _01067_ _01057_ _00611_ VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__mux2_1
X_09735_ _03633_ _03641_ _03642_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__o21ai_1
X_09666_ H\[2\]\[6\] _03022_ _03574_ VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06878_ result_reg_Rshift\[11\] _00753_ _01001_ VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__o21ai_1
X_08617_ _02523_ Qset\[0\]\[0\] VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _03505_ VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_25_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _02462_ _02465_ VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__nand2_1
X_08479_ H\[1\]\[10\] VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__inv_2
X_11490_ _05380_ _05390_ VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__or2_1
X_10510_ H\[3\]\[9\] _03792_ _03794_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_33_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10441_ _03652_ _03868_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10372_ _04203_ _04264_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__nor2_1
X_12111_ result_reg_and\[8\] _05894_ _05920_ _05921_ _02125_ VGND VGND VPWR VPWR _00348_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12042_ result_reg_Rshift\[12\] _05847_ VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_5_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12944_ clknet_leaf_21_clk _00387_ VGND VGND VPWR VPWR result_reg_not\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_130 _05717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12875_ clknet_leaf_24_clk _00318_ VGND VGND VPWR VPWR result_reg_Lshift\[10\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_141 _06284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_152 R2\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_163 _00396_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_174 _01670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11826_ result_reg_mul\[13\] _05669_ _05682_ VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__o21ai_1
XANTENNA_185 im_reg\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11757_ _05628_ _04256_ _05647_ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10708_ H\[3\]\[10\] _03792_ _03794_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11688_ _05572_ _05587_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10639_ _02567_ _02384_ VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12309_ result_reg_set\[7\] _06063_ _06066_ _06072_ VGND VGND VPWR VPWR _00395_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07850_ result_reg_mul\[14\] _01679_ _01656_ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__o21ai_1
X_07781_ _01716_ _00975_ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__nand2_1
X_06801_ _00927_ Qset\[0\]\[8\] _00687_ VGND VGND VPWR VPWR _00928_ sky130_fd_sc_hd__mux2_1
Xinput3 data_in[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
X_06732_ _00860_ _00745_ VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__or2_1
X_09520_ _03426_ _03427_ _03026_ _03428_ _03429_ VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__a32o_1
XFILLER_0_78_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06663_ net11 _00696_ _00793_ VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__o21ai_1
X_09451_ _03359_ _03360_ VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__nand2_1
X_06594_ result_reg_mul\[2\] VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__inv_2
X_09382_ _03291_ _03292_ VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__nor2_2
X_08402_ _02322_ _02325_ VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08333_ _02230_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__buf_6
X_08264_ _02193_ net55 _02170_ VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07215_ result_reg_Lshift\[3\] result_reg_Rshift\[3\] _01165_ VGND VGND VPWR VPWR
+ _01297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08195_ _00591_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_30_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07146_ _00557_ _00631_ _01230_ VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07077_ _01157_ VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07979_ Oset\[0\]\[0\] _01218_ _02001_ VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__mux2_1
X_09718_ _03619_ _03624_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__nand2_1
X_10990_ _00498_ _00585_ _04887_ _04892_ _03768_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_2_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09649_ _03553_ VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12660_ clknet_leaf_53_clk _00110_ VGND VGND VPWR VPWR Oset\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_11611_ _05335_ H\[1\]\[15\] VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12591_ clknet_leaf_46_clk _00041_ VGND VGND VPWR VPWR Qset\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11542_ _05442_ VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__inv_2
X_11473_ _05360_ _05373_ VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__or2_1
X_10424_ _04329_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10355_ _04199_ _04221_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10286_ _04159_ _04192_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__or2_1
X_12025_ _05855_ VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12927_ clknet_leaf_30_clk _00370_ VGND VGND VPWR VPWR result_reg_or\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12858_ clknet_leaf_18_clk _00301_ VGND VGND VPWR VPWR result_reg_mac\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11809_ result_reg_mul\[7\] _05669_ _05682_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12789_ clknet_leaf_53_clk _00232_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07000_ _01114_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08951_ _02737_ _02829_ VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__nor2_1
X_08882_ _00681_ _00580_ _02539_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__o21ai_1
X_07902_ Oset\[2\]\[4\] _01332_ _01942_ VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__mux2_1
X_07833_ net5 _01746_ VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_16_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07764_ _01819_ H\[3\]\[9\] _01629_ VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07695_ result_reg_or\[6\] _01595_ VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__nor2_1
X_06715_ _00844_ _00735_ VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__nand2_1
X_09503_ _03379_ _00623_ _03412_ VGND VGND VPWR VPWR _03413_ sky130_fd_sc_hd__nand3_1
X_06646_ result_reg_not\[3\] VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09434_ H\[2\]\[5\] H\[3\]\[5\] _02611_ VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06577_ _00662_ CMD_and _00527_ VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__or3_1
X_09365_ _03273_ _03274_ _03275_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__nand3_1
XANTENNA_41 _01059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_30 _00878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Left_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08316_ _02240_ _02143_ _02242_ VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__nand3_1
X_09296_ _03205_ _03206_ VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_74 _01502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 _01410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 _01278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08247_ _02175_ _02135_ _02176_ VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__nand3_1
XFILLER_0_34_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_96 _01811_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 _01731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08178_ _02102_ _02103_ net46 VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_76_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07129_ _01213_ VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__clkbuf_4
X_10140_ _04042_ _04043_ _04044_ _04046_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__a2bb2o_2
XTAP_TAPCELL_ROW_7_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10071_ _03972_ _03973_ _03977_ VGND VGND VPWR VPWR _03978_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_34_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10973_ _04830_ _04854_ _04875_ VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12712_ clknet_leaf_52_clk _00155_ VGND VGND VPWR VPWR Oset\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12643_ clknet_leaf_51_clk _00093_ VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_53_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12574_ clknet_leaf_49_clk _00024_ VGND VGND VPWR VPWR Qset\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11525_ _05424_ _05425_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11456_ _04830_ _05341_ _05356_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11387_ _05287_ _05288_ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10407_ _04263_ _04311_ _04312_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__nand3b_1
X_10338_ _04242_ _04243_ _04244_ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__nand3_1
X_12008_ _00640_ _05667_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__nand2_2
X_10269_ _04147_ _04175_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07480_ _01544_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__clkbuf_4
X_06500_ _00634_ VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__buf_4
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06431_ _00565_ VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09150_ _02561_ _02323_ VGND VGND VPWR VPWR _03061_ sky130_fd_sc_hd__nor2_1
X_06362_ _00495_ _00500_ VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__nand2_1
X_06293_ _06259_ net64 VGND VGND VPWR VPWR _06260_ sky130_fd_sc_hd__nand2_1
X_08101_ _01819_ H\[1\]\[9\] _02057_ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__mux2_1
X_09081_ _02586_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__buf_6
X_08032_ _02029_ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09983_ _03877_ _03889_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08934_ Qset\[2\]\[2\] Qset\[3\]\[2\] _02625_ VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__mux2_1
X_08865_ _02586_ H\[3\]\[2\] _02591_ _02777_ VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07816_ result_reg_mul\[12\] _01585_ _01589_ VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__o21ai_1
X_08796_ _02708_ _02533_ _02709_ VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__nand3_1
X_07747_ result_reg_mac\[9\] _01541_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07678_ result_reg_Rshift\[5\] _01672_ _01607_ _01737_ VGND VGND VPWR VPWR _01738_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06629_ result_reg_mac\[3\] VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09417_ _03325_ _02991_ _03326_ VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__nand3_1
X_09348_ _03205_ _03258_ VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11310_ _04494_ _04982_ _04690_ _04957_ VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_10_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09279_ _03116_ _03106_ VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12290_ _06058_ R2\[0\] VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11241_ _04832_ Qset\[2\]\[13\] VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__nor2_1
X_11172_ _05073_ _05072_ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__nand2_1
X_10123_ _04028_ _04029_ VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_89_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10054_ _03957_ _03960_ VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_46_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10956_ _03795_ VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10887_ _04788_ _04790_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12626_ clknet_leaf_45_clk _00076_ VGND VGND VPWR VPWR Oset\[3\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12557_ _06249_ VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__clkbuf_1
X_12488_ _01147_ _05134_ VGND VGND VPWR VPWR _06210_ sky130_fd_sc_hd__and2_1
X_11508_ _05358_ _05408_ VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__nand2_1
X_11439_ _05333_ _03758_ _00589_ _05339_ VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06980_ _01082_ _00695_ _01091_ _01099_ _00644_ VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__a221o_1
X_08650_ _02562_ VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__buf_4
X_07601_ result_reg_mul\[2\] _01663_ _01589_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08581_ _02311_ _02482_ _02139_ _02489_ _02497_ VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_44_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07532_ _01574_ _01592_ _01594_ _01596_ VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_105_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07463_ _01530_ VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_105_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06414_ _00548_ VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__buf_4
X_09202_ _03111_ _03112_ VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__nand2_1
X_07394_ _01010_ _01466_ _01177_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__mux2_1
X_09133_ _01537_ _03043_ VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__nor2_1
X_06345_ R2\[0\] _00486_ VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09064_ Oset\[1\]\[3\] _02836_ VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08015_ Oset\[1\]\[1\] _01278_ _02019_ VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09966_ _02396_ _02544_ VGND VGND VPWR VPWR _03873_ sky130_fd_sc_hd__nand2_1
X_08917_ _02829_ _02737_ VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__nand2_1
X_09897_ _03801_ _03794_ _00647_ _03803_ VGND VGND VPWR VPWR _03804_ sky130_fd_sc_hd__a211o_1
X_08848_ _02760_ _00580_ VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08779_ Qset\[2\]\[1\] Qset\[3\]\[1\] _02624_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _01148_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_43_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _04711_ _04713_ VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10741_ _04517_ _04521_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12411_ _06149_ net23 _06139_ VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__a21o_1
X_10672_ _03350_ _04050_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_20_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_51_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12342_ _06092_ VGND VGND VPWR VPWR _00408_ sky130_fd_sc_hd__clkbuf_1
X_12273_ _06032_ _01024_ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11224_ _05122_ _05126_ _04816_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__nand3_1
X_11155_ _05056_ _05057_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11086_ _04979_ _04988_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__or2_1
X_10106_ _03505_ _03876_ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__nand2_1
X_10037_ _03941_ _03943_ VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_59_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11988_ _04963_ _00590_ _04047_ _05749_ _05826_ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10939_ _04837_ _04839_ _03764_ _04840_ _04841_ VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_11_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12609_ clknet_leaf_48_clk _00059_ VGND VGND VPWR VPWR Qset\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09820_ _03727_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__inv_2
X_06963_ result_reg_add\[15\] VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__inv_2
X_09751_ _03655_ _03658_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__nand2_1
X_08702_ _02610_ _02616_ VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__nand2_1
X_06894_ _01016_ _01007_ _00730_ VGND VGND VPWR VPWR _01017_ sky130_fd_sc_hd__mux2_1
X_09682_ _00623_ _03506_ _03590_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_55_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08633_ Oset\[1\]\[0\] _02529_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__nand2_1
X_08564_ _02459_ Qset\[1\]\[14\] _02444_ _02480_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07515_ _01579_ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08495_ _02364_ Oset\[3\]\[11\] _02347_ _02414_ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__a211o_1
X_07446_ _01512_ _01515_ _01271_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07377_ _01450_ _01187_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06328_ _00472_ current_state\[6\] VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__nand2_2
XFILLER_0_44_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09116_ _03026_ VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09047_ _00549_ _02957_ _02958_ VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09949_ _03849_ _03855_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12960_ clknet_leaf_2_clk _00403_ VGND VGND VPWR VPWR result_reg_set\[15\] sky130_fd_sc_hd__dfxtp_1
X_12891_ clknet_leaf_24_clk _00334_ VGND VGND VPWR VPWR result_reg_Rshift\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_28_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ _02866_ _02869_ VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__nand2_1
X_11842_ _05706_ _02750_ VGND VGND VPWR VPWR _05708_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_56_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11773_ _05315_ _05316_ _05655_ _05658_ VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10724_ _01537_ _04614_ _04616_ _00556_ _04628_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__a311o_2
XFILLER_0_82_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10655_ _04539_ _04559_ VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12325_ result_reg_set\[13\] _06063_ _06066_ _06082_ VGND VGND VPWR VPWR _00401_
+ sky130_fd_sc_hd__o211a_1
X_10586_ _03758_ _04490_ VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12256_ _06032_ _05769_ _06013_ _06038_ VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12187_ _05937_ _05909_ _05984_ _05957_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__a211o_1
X_11207_ _05108_ _05109_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__nand2_1
X_11138_ _05040_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__inv_2
X_11069_ _04048_ _03745_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_0_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07300_ _01267_ _00883_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08280_ _02151_ _02207_ _02147_ _02208_ VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__a211o_1
X_07231_ _00761_ _01275_ _01276_ VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07162_ _00567_ _01243_ _01220_ _01245_ _01246_ VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07093_ _00609_ _01175_ _01177_ VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09803_ H\[2\]\[7\] _03023_ _03710_ VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__a21o_1
X_07995_ Oset\[0\]\[8\] _01403_ _02001_ VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__mux2_1
X_06946_ result_reg_sub\[14\] VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__inv_2
X_09734_ _02326_ _00584_ _02573_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__a21oi_1
X_06877_ _00754_ _01000_ VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09665_ H\[3\]\[6\] _03033_ _03026_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__a21o_1
X_08616_ _02524_ _02526_ _02530_ VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__nand3_1
XFILLER_0_77_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ _03504_ _02308_ VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_25_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _02459_ Oset\[1\]\[13\] _02378_ _02464_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__a211o_1
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08478_ _02396_ _02373_ _02374_ _02398_ VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__a211o_1
X_07429_ result_reg_add\[14\] _01202_ VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10440_ _04345_ _04025_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10371_ _04203_ _04264_ _04276_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12110_ _05881_ _03824_ _03775_ _05894_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_20_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12041_ _05864_ VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12943_ clknet_leaf_26_clk _00386_ VGND VGND VPWR VPWR result_reg_not\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_5_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 _05721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12874_ clknet_leaf_24_clk _00317_ VGND VGND VPWR VPWR result_reg_Lshift\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_120 _03449_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_142 _06284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_175 _01771_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_164 _00414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11825_ _05695_ VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__inv_2
XANTENNA_153 R2\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11756_ _05628_ _00912_ _02650_ VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_186 _00809_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10707_ _04610_ _04611_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__nand2_1
X_11687_ _05585_ _05586_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__xor2_1
XFILLER_0_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10638_ _04542_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__inv_2
X_10569_ _04282_ Qset\[3\]\[10\] _03761_ _04473_ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__a211o_1
X_12308_ _06058_ _06071_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12239_ _05958_ _06026_ VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__nand2_1
X_07780_ _01834_ result_reg_mac\[10\] _01570_ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__mux2_1
X_06800_ _00918_ _00645_ _00920_ _00926_ VGND VGND VPWR VPWR _00927_ sky130_fd_sc_hd__a31o_4
Xinput4 data_in[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
X_06731_ result_reg_mul\[6\] VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09450_ _03357_ _03352_ _03353_ VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__nand3_1
XFILLER_0_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06662_ _00792_ _00735_ VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__nand2_1
X_08401_ _02319_ Oset\[1\]\[7\] _02250_ _02324_ VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__a211o_1
X_06593_ result_reg_set\[2\] VGND VGND VPWR VPWR _00726_ sky130_fd_sc_hd__inv_2
X_09381_ _03290_ _03046_ VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08332_ _02258_ _02250_ VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08263_ _02126_ _02178_ _02140_ _02185_ _02192_ VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_46_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07214_ _01296_ VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08194_ net37 _02124_ _02125_ VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07145_ shift.left CMD_logic_shift_right _00624_ _01229_ VGND VGND VPWR VPWR _01230_
+ sky130_fd_sc_hd__or4_1
XFILLER_0_6_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07076_ _01160_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_98_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07978_ _02000_ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__buf_4
X_06929_ _00754_ _01050_ VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__nand2_1
X_09717_ _03611_ _03619_ _03624_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09648_ _03553_ _03555_ _03556_ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_38_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _03001_ _02289_ _02991_ _03487_ VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__o211ai_1
X_11610_ _05335_ _02514_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__nor2_1
X_12590_ clknet_leaf_49_clk _00040_ VGND VGND VPWR VPWR Qset\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_11541_ _05440_ _05441_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11472_ _05371_ _05372_ VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10423_ _03859_ _02620_ _03745_ _03835_ _03908_ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__a32o_1
XFILLER_0_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10354_ _04244_ _04239_ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__nand2_1
X_10285_ _04190_ _04191_ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12024_ _00805_ _05844_ _05775_ _05854_ VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__a211o_1
X_12926_ clknet_leaf_16_clk _00369_ VGND VGND VPWR VPWR result_reg_or\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ clknet_leaf_10_clk _00300_ VGND VGND VPWR VPWR result_reg_mac\[8\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11808_ _05684_ VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12788_ clknet_leaf_54_clk _00231_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11739_ _00728_ _05628_ _05634_ _05635_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__a211o_1
XFILLER_0_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08950_ _02862_ VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__inv_2
X_07901_ _01946_ VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__clkbuf_1
X_08881_ _02790_ _02793_ _00581_ VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__nand3_1
X_07832_ _01033_ _01682_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__or2_1
X_07763_ _01803_ _01815_ _01613_ _01818_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_79_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09502_ _03411_ _03233_ VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__nand2_1
X_07694_ _01691_ result_reg_and\[6\] VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__nand2_1
X_06714_ _00840_ _00843_ _00608_ VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06645_ _00761_ _00695_ _00776_ _00725_ _00644_ VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__a221o_1
X_09433_ H\[1\]\[5\] _03341_ _02591_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__o21a_1
X_09364_ _03267_ _03272_ _03271_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__nand3_1
X_06576_ _00624_ VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__buf_6
X_08315_ _02241_ Qset\[3\]\[4\] VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_20 _00759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 _00904_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09295_ _03176_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_53 _01284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 _01432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_75 _01507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_42 _01072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08246_ _02127_ Qset\[1\]\[1\] VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__nand2_1
XANTENNA_86 _01744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08177_ im_reg\[7\] _02100_ _02105_ _02112_ VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__o211a_1
XANTENNA_97 _01819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07128_ _00647_ _00625_ _00627_ VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_76_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07059_ current_state\[2\] VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_7_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10070_ _03975_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10972_ _01538_ _04861_ _04864_ _02096_ _04874_ VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__a311o_2
XFILLER_0_97_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12711_ clknet_leaf_45_clk _00154_ VGND VGND VPWR VPWR Oset\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_12642_ clknet_leaf_51_clk _00092_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12573_ clknet_leaf_28_clk _00023_ VGND VGND VPWR VPWR next_PC\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11524_ _04895_ _05379_ _05423_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_13_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11455_ _01538_ _05343_ _05345_ _02096_ _05355_ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__a311o_2
XFILLER_0_68_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10406_ _04310_ _04277_ _04279_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_33_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11386_ _05286_ _05284_ VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__nand2_1
X_10337_ _04241_ _04240_ VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10268_ _04173_ _04174_ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__nand2_1
X_12007_ _05774_ _05841_ _05808_ _05842_ VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__o211a_1
X_10199_ _04105_ H\[3\]\[12\] _04045_ VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12909_ clknet_leaf_31_clk _00352_ VGND VGND VPWR VPWR result_reg_and\[12\] sky130_fd_sc_hd__dfxtp_2
X_06430_ _00471_ CMD_addition current_state\[5\] VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06361_ _00500_ _00495_ VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__or2_1
X_06292_ net35 VGND VGND VPWR VPWR _06259_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08100_ _02066_ VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__clkbuf_1
X_09080_ _02584_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__buf_4
X_08031_ Oset\[1\]\[9\] _01420_ _02019_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09982_ _02619_ _03868_ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__nand2_1
X_08933_ _02837_ _02843_ _02845_ VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08864_ _02592_ _02207_ VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__nor2_1
X_07815_ _01586_ result_reg_sub\[12\] VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__nand2_1
X_08795_ _02527_ Qset\[1\]\[1\] VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07746_ _01802_ VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07677_ _01716_ _00850_ VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__nand2_1
X_09416_ _02992_ Qset\[3\]\[5\] VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06628_ _00760_ VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__clkbuf_1
X_06559_ _00689_ _00692_ _00656_ VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__mux2_1
X_09347_ _03257_ VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09278_ _03183_ _03186_ _03188_ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08229_ _02092_ VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_10_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11240_ _03770_ _05141_ _01156_ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__o21ai_1
X_11171_ _05072_ _05073_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__or2_1
X_10122_ _04027_ _04011_ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10053_ _03958_ _03919_ _03959_ VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10955_ _04857_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10886_ _04789_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12625_ clknet_leaf_45_clk _00075_ VGND VGND VPWR VPWR Oset\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12556_ _01080_ Qset\[3\]\[14\] _06233_ VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__mux2_1
X_11507_ _05407_ VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__inv_2
X_12487_ _06209_ _06202_ VGND VGND VPWR VPWR _00436_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11438_ _03758_ _05338_ VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__nor2_1
X_11369_ _05256_ _05270_ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07600_ _01584_ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__clkbuf_4
X_08580_ _02493_ _02496_ _01554_ VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__a21o_2
XPHY_EDGE_ROW_53_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07531_ result_reg_or\[0\] _01595_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07462_ _01529_ _01149_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07393_ _01016_ _01007_ _01174_ VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__mux2_1
X_06413_ CMD_mul_accumulation VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__inv_2
X_09201_ _03080_ _03076_ VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06344_ _00484_ _00485_ _00486_ VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__a21bo_1
X_09132_ _03037_ _03042_ _00621_ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_62_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09063_ _02632_ Oset\[0\]\[3\] _02840_ VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08014_ _02020_ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09965_ _02561_ H\[2\]\[10\] _02727_ VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__o21a_1
X_09896_ Oset\[3\]\[8\] _03023_ _03798_ _03802_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__o211a_1
X_08916_ _02786_ _02825_ VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_71_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08847_ _02756_ _02759_ VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__nand2_2
XFILLER_0_79_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08778_ H\[1\]\[1\] _02688_ _00001_ _02691_ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__a211o_1
X_07729_ _01390_ _01682_ VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10740_ _04644_ VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_84_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10671_ _04124_ _04369_ _04372_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__o21a_1
X_12410_ _06128_ _06116_ VGND VGND VPWR VPWR _06149_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_80_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12341_ _06091_ _01532_ VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__and2_1
X_12272_ _06039_ _05817_ _06044_ _06047_ VGND VGND VPWR VPWR _00383_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_95_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11223_ _05123_ _05124_ _05125_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11154_ _04175_ _04147_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__nand2_1
X_10105_ _03994_ _03990_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__and2_1
X_11085_ _04986_ _04987_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__nand2_1
X_10036_ _03942_ _03923_ VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_59_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11987_ _01162_ _05825_ VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10938_ _03773_ _02439_ VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10869_ _04771_ _04772_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__and2b_1
X_12608_ clknet_leaf_46_clk _00058_ VGND VGND VPWR VPWR Qset\[2\]\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_5_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12539_ _06240_ VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06962_ result_reg_mac\[15\] VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__inv_2
X_09750_ _03656_ _03657_ _03653_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__nand3_1
XFILLER_0_39_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09681_ _01537_ _03575_ _03577_ _00549_ _03589_ VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__a311o_2
X_08701_ _02613_ _02615_ _02571_ VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__nand3_1
X_06893_ result_reg_sub\[12\] VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08632_ _02545_ _02142_ _02526_ _02546_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__o211ai_1
X_08563_ _02459_ _02479_ VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__nor2_1
X_07514_ _01578_ _00537_ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__nor2_4
XFILLER_0_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08494_ _02356_ _02413_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__nor2_1
X_07445_ _01086_ _01266_ _01299_ _01514_ VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07376_ _01447_ _01449_ _01182_ VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__mux2_1
X_06327_ _00471_ VGND VGND VPWR VPWR _00472_ sky130_fd_sc_hd__buf_2
X_09115_ _02837_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__buf_2
XFILLER_0_17_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09046_ _02895_ _00549_ VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09948_ _03854_ _02573_ _00588_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09879_ _00584_ _03785_ VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__nor2_1
X_12890_ clknet_leaf_23_clk _00333_ VGND VGND VPWR VPWR result_reg_Rshift\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11910_ _05744_ _02711_ _05758_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__a21o_2
X_11841_ _05706_ VGND VGND VPWR VPWR _05707_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_56_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _05627_ _01035_ _02115_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__a21o_1
X_10723_ _01537_ _04627_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10654_ _04557_ _04558_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__nor2b_1
XTAP_TAPCELL_ROW_97_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10585_ _03764_ _04487_ _04488_ _04489_ VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__o2bb2a_1
X_12324_ R1\[1\] _05745_ R3\[1\] _05744_ _06054_ VGND VGND VPWR VPWR _06082_ sky130_fd_sc_hd__a221o_1
X_12255_ _06033_ _00804_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12186_ _05888_ _03346_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__nor2_1
X_11206_ _05107_ _05060_ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__nand2_1
X_11137_ _05038_ _05039_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__nand2_1
X_11068_ _04964_ _01156_ _04970_ _03132_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__a31o_1
X_10019_ _03883_ _03878_ VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07230_ _01192_ _01304_ _01305_ _01275_ _01311_ VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__a311o_1
XFILLER_0_41_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07161_ _01159_ _01202_ _01208_ _01190_ VGND VGND VPWR VPWR _01246_ sky130_fd_sc_hd__or4_1
XFILLER_0_54_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07092_ _01176_ VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__buf_4
XFILLER_0_41_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09802_ H\[3\]\[7\] _03025_ _03027_ VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__a21o_1
X_07994_ _02009_ VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__clkbuf_1
X_06945_ result_reg_set\[14\] VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__inv_2
X_09733_ _03634_ _03640_ _02540_ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__and3_1
X_06876_ result_reg_Lshift\[11\] VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__inv_2
X_09664_ _03571_ _00831_ _03572_ VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__nand3_1
XFILLER_0_96_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09595_ _03496_ _03503_ VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__nand2_2
X_08615_ Qset\[3\]\[0\] _02529_ VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ _02459_ _02463_ VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08477_ _02397_ H\[2\]\[10\] VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07428_ result_reg_and\[14\] VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07359_ _01433_ _01238_ _01215_ VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10370_ _04272_ _04275_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_79_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09029_ _02592_ _02234_ VGND VGND VPWR VPWR _02941_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_92_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12040_ _05822_ _05851_ _05775_ _05863_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__a211o_1
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12942_ clknet_leaf_26_clk _00385_ VGND VGND VPWR VPWR result_reg_not\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_121 _03601_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_132 _05725_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12873_ clknet_leaf_24_clk _00316_ VGND VGND VPWR VPWR result_reg_Lshift\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_110 _02116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_143 _06284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_176 _01785_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11824_ _05054_ _05115_ _05677_ _05694_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__a31o_1
XANTENNA_165 _00498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_154 R2\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11755_ _05646_ VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_187 _00809_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10706_ _04606_ _02092_ _04608_ VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__nand3_1
X_11686_ _05397_ _05394_ _05395_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__a21bo_1
X_10637_ _02567_ Oset\[1\]\[10\] VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__nand2_1
X_10568_ _03759_ _04472_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12307_ _00671_ _02311_ _01990_ _02139_ _03075_ VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__o221a_1
X_10499_ _03859_ _02096_ VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__nand2_1
X_12238_ _05500_ _04086_ _05881_ VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__a21o_1
X_12169_ _02807_ _05889_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__nand2_1
Xinput5 data_in[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
X_06730_ result_reg_sub\[6\] _00541_ _00858_ VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__o21ai_1
X_06661_ _00786_ _00791_ _00608_ VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__mux2_1
X_08400_ _02261_ _02323_ VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06592_ _00628_ VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__clkbuf_4
X_09380_ _03046_ _03290_ VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__nor2_4
X_08331_ H\[2\]\[4\] H\[3\]\[4\] _02241_ VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__mux2_1
X_08262_ _02188_ _02191_ _01551_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__a21o_1
X_07213_ Oset\[3\]\[2\] _01295_ _01250_ VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__mux2_1
X_08193_ _01148_ VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__buf_4
XFILLER_0_54_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07144_ CMD_not _00545_ CMD_and _01228_ VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__or4_1
X_07075_ _01159_ VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__buf_2
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07977_ _01940_ _01999_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__nor2_4
X_06928_ result_reg_Lshift\[13\] VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__inv_2
X_09716_ _03621_ _03622_ _03623_ VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__nand3_2
XFILLER_0_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06859_ _00740_ _00982_ _00535_ VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__a21oi_1
X_09647_ _03395_ _03394_ _03401_ VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_38_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09578_ _03001_ Qset\[3\]\[6\] VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__nand2_1
X_08529_ _02446_ _02373_ _02378_ _02447_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__a211o_1
XFILLER_0_65_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11540_ _03051_ _04607_ _04924_ VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__or3_1
XFILLER_0_25_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11471_ _05370_ _05361_ VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__nand2_1
X_10422_ _04325_ _04327_ VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__nand2_1
X_10353_ _04259_ VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12023_ _05844_ _05780_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__nor2_1
X_10284_ _04185_ _04183_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__or2_1
X_12925_ clknet_leaf_21_clk _00368_ VGND VGND VPWR VPWR result_reg_or\[12\] sky130_fd_sc_hd__dfxtp_1
X_12856_ clknet_leaf_18_clk _00299_ VGND VGND VPWR VPWR result_reg_mac\[7\] sky130_fd_sc_hd__dfxtp_1
X_11807_ _03569_ _03570_ _05677_ _05683_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12787_ clknet_leaf_54_clk _00230_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dfxtp_1
X_11738_ _05631_ _02860_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11669_ _05560_ _05568_ VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08880_ _02791_ _02535_ _02792_ VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__nand3_2
X_07900_ Oset\[2\]\[3\] _01314_ _01942_ VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__mux2_1
X_07831_ _01881_ _01653_ _01882_ VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07762_ _00948_ _01607_ _01817_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__o21ai_1
X_09501_ _03407_ _03410_ VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__nand2_2
X_07693_ _01749_ _01663_ _01750_ _01751_ VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__a31o_1
X_06713_ _00815_ _00842_ _00613_ VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06644_ _00739_ _00768_ _00769_ _00774_ _00775_ VGND VGND VPWR VPWR _00776_ sky130_fd_sc_hd__a32o_1
X_09432_ _03341_ _02281_ VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_35_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06575_ _00552_ VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__buf_2
XFILLER_0_59_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09363_ _03079_ VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08314_ _02131_ VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__buf_6
XANTENNA_21 _00776_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 _00649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_32 _00904_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09294_ _03020_ VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_54 _01325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 _01074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08245_ _02128_ Qset\[0\]\[1\] VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__nand2_1
XANTENNA_65 _01437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_87 _01752_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 _01565_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08176_ _02102_ _02103_ net45 VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__a21o_1
XANTENNA_98 _01819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07127_ result_reg_or\[0\] _01199_ _01192_ _01211_ VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07058_ _01145_ VGND VGND VPWR VPWR _00071_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10971_ _04868_ _04873_ _01538_ VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_87_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12710_ clknet_leaf_53_clk _00153_ VGND VGND VPWR VPWR Oset\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_12641_ clknet_leaf_52_clk _00091_ VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_65_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12572_ clknet_leaf_34_clk _00022_ VGND VGND VPWR VPWR next_PC\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11523_ _04895_ _05379_ _05423_ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_41_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11454_ _05349_ _05354_ _01538_ VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__a21oi_1
X_10405_ _04280_ _04310_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11385_ _05284_ _05286_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__or2_1
X_10336_ _03949_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10267_ _03922_ _03956_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__nand2_1
X_12006_ _05774_ _01103_ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__nand2_1
X_10198_ _02567_ VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_49_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12908_ clknet_leaf_16_clk _00351_ VGND VGND VPWR VPWR result_reg_and\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12839_ clknet_leaf_0_clk _00282_ VGND VGND VPWR VPWR result_reg_mul\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_33_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06360_ next_PC\[5\] VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__inv_2
X_06291_ _06253_ _06254_ _06257_ VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__or3_2
X_08030_ _02028_ VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput30 instruction_in[5] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_1
XFILLER_0_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09981_ _03880_ _03887_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__or2_1
X_08932_ Oset\[0\]\[2\] _02632_ _02844_ VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__a21o_1
X_08863_ _02775_ _02555_ VGND VGND VPWR VPWR _02776_ sky130_fd_sc_hd__nand2_1
X_07814_ _01581_ result_reg_add\[12\] VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08794_ _02522_ Qset\[0\]\[1\] VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__nand2_1
X_07745_ _01801_ H\[3\]\[8\] _01629_ VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__mux2_1
X_07676_ _01735_ result_reg_mac\[5\] _01570_ VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__mux2_1
X_09415_ _02582_ Qset\[2\]\[5\] VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06627_ _00759_ Qset\[0\]\[2\] _00687_ VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__mux2_1
X_06558_ _00690_ _00691_ _00643_ VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09346_ _03051_ _02578_ VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__nor2_1
X_06489_ _00623_ VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__buf_4
X_09277_ _03187_ VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__inv_2
X_08228_ _02126_ _02138_ _02140_ _02150_ _02158_ VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__o221ai_4
X_08159_ _02095_ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__buf_2
X_11170_ _03383_ _03507_ _03692_ _03689_ VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__o31a_1
XFILLER_0_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10121_ _04011_ _04027_ VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__or2_1
X_10052_ _03924_ _03942_ VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_89_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10954_ _03793_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__clkbuf_4
X_10885_ _04759_ _04760_ _03751_ _03745_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__a31o_1
X_12624_ clknet_leaf_53_clk _00074_ VGND VGND VPWR VPWR Oset\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12555_ _06248_ VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11506_ _05405_ _05406_ VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12486_ _06102_ Qim _04827_ VGND VGND VPWR VPWR _06209_ sky130_fd_sc_hd__o21ai_1
X_11437_ _05334_ _05336_ _05337_ _04835_ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11368_ _05257_ _05269_ VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10319_ _03666_ _03518_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__nand2_1
X_11299_ _05199_ _05195_ _05196_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_28_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07530_ _01572_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07461_ R2\[1\] net28 current_state\[2\] VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__mux2_1
X_07392_ result_reg_set\[12\] VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__inv_2
X_06412_ CMD_and VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__inv_2
X_09200_ _03052_ _03110_ VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06343_ _06284_ VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__buf_2
XFILLER_0_44_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09131_ _03038_ _03039_ _03027_ _03040_ _03041_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__a32o_1
XFILLER_0_44_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09062_ _02632_ Oset\[2\]\[3\] VGND VGND VPWR VPWR _02974_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08013_ Oset\[1\]\[0\] _01218_ _02019_ VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09964_ _02400_ _02874_ VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__nand2_1
X_09895_ Oset\[2\]\[8\] _03791_ VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__or2_1
X_08915_ _02737_ _02826_ _02827_ VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__nand3b_2
X_08846_ _02757_ _02590_ _02758_ VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__nand3_1
X_08777_ _02688_ _02189_ VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__nor2_1
X_07728_ _01783_ _01653_ _01784_ VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__a21o_1
X_07659_ _01715_ _01719_ _01613_ VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_84_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10670_ _03507_ _04110_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09329_ _02783_ _02213_ _02897_ VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_51_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12340_ im_reg\[7\] net32 _01146_ VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__mux2_1
X_12271_ _06032_ _00999_ VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11222_ _04633_ _04820_ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__nor2_1
X_11153_ _04176_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__inv_2
X_11084_ _04495_ _04975_ _04985_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__o21ai_1
X_10104_ _04002_ _03997_ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__and2_1
X_10035_ _03940_ _03938_ VGND VGND VPWR VPWR _03942_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_59_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11986_ _04969_ VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10937_ Oset\[1\]\[12\] _03773_ _03761_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12607_ clknet_leaf_46_clk _00057_ VGND VGND VPWR VPWR Qset\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_10868_ _04770_ _04764_ VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10799_ _04697_ _04699_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12538_ _00854_ Qset\[3\]\[5\] _06234_ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__mux2_1
X_12469_ _06097_ Oreg2 _06195_ _06197_ _02101_ VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__o221a_1
XFILLER_0_41_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06961_ _01081_ VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__clkbuf_1
X_09680_ _01536_ _03588_ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__nor2_1
X_08700_ _02586_ H\[1\]\[0\] _02584_ _02614_ VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__a211o_1
X_06892_ _01014_ _00553_ VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__or2_1
X_08631_ Oset\[3\]\[0\] _02545_ VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08562_ Qset\[0\]\[14\] VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__inv_2
X_07513_ _01571_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__clkinv_4
X_08493_ Oset\[2\]\[11\] VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__inv_2
X_07444_ _01093_ _01267_ _01263_ _01513_ VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07375_ _00985_ _01448_ _01177_ VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06326_ _06259_ _06263_ _06271_ VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__and3_2
X_09114_ _03024_ VGND VGND VPWR VPWR _03025_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09045_ _02954_ _02956_ VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09947_ _02560_ _03850_ _03851_ _03853_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__o31a_2
XFILLER_0_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09878_ _03770_ _03775_ _03784_ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08829_ _00536_ _02742_ VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__xor2_1
X_11840_ _05702_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _05657_ VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10722_ _04621_ _04626_ _00621_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10653_ _04556_ _04347_ VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__nand2_1
X_10584_ H\[1\]\[10\] _04302_ _03761_ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12323_ result_reg_set\[12\] _06063_ _06066_ _06081_ VGND VGND VPWR VPWR _00400_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12254_ _05762_ _06033_ _06013_ _06037_ VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12185_ _05881_ _03122_ _05888_ _03141_ _05982_ VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__o221ai_1
X_11205_ _05060_ _05107_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__or2_1
X_11136_ _05037_ _05036_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__nand2_1
X_11067_ _04969_ _03781_ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__nand2_1
X_10018_ _03897_ _03350_ _03898_ VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__or3_1
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11969_ _00590_ _04552_ _04546_ _01158_ _05810_ VGND VGND VPWR VPWR _05811_ sky130_fd_sc_hd__a221oi_4
XTAP_TAPCELL_ROW_102_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07160_ _01244_ VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__buf_4
XFILLER_0_6_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07091_ _01172_ _00532_ VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__nand2_4
XFILLER_0_14_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09801_ _03705_ _02092_ _03706_ VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__nand3_1
XFILLER_0_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07993_ Oset\[0\]\[7\] _01385_ _02001_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__mux2_1
X_09732_ _03639_ _00581_ VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__nand2_1
X_06944_ _01063_ _01064_ _00835_ VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__a21o_1
X_06875_ result_reg_not\[11\] VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__inv_2
X_09663_ _00623_ _03110_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08614_ _02528_ VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__buf_6
X_09594_ _03502_ _02573_ _00587_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__a21oi_1
X_08545_ Oset\[0\]\[13\] VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_53_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08476_ _02356_ VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__buf_4
XFILLER_0_92_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07427_ _01496_ _01193_ _01191_ _01497_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__a211o_1
XFILLER_0_64_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07358_ _01429_ _01432_ _00965_ _01271_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_45_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06309_ current_state\[4\] VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07289_ _01161_ _01352_ _01367_ VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__a21bo_4
XFILLER_0_32_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09028_ _02592_ H\[3\]\[3\] _02591_ _02939_ VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__a211o_1
XFILLER_0_32_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12941_ clknet_leaf_26_clk _00384_ VGND VGND VPWR VPWR result_reg_not\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ clknet_leaf_22_clk _00315_ VGND VGND VPWR VPWR result_reg_Lshift\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_100 _01823_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_122 _03601_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_133 _05792_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11823_ result_reg_mul\[12\] _05669_ _05682_ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__o21ai_1
XANTENNA_111 _02168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_166 _00498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_144 im_reg\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_155 R2\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11754_ _00883_ _05631_ _05634_ _05645_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__a211o_1
XANTENNA_177 _01883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_188 _00809_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10705_ _04609_ _00831_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__nand2_1
X_11685_ _05573_ _05584_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__xor2_1
XFILLER_0_102_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10636_ _04105_ _02387_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10567_ Qset\[2\]\[10\] VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__inv_2
X_12306_ result_reg_set\[6\] _06063_ _06066_ _06070_ VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__o211a_1
X_10498_ _04338_ _00710_ _04403_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__nand3_1
X_12237_ result_reg_or\[14\] _05960_ _06023_ _06025_ _02101_ VGND VGND VPWR VPWR _00370_
+ sky130_fd_sc_hd__o221a_1
X_12168_ _05750_ _02760_ _05907_ VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__a21oi_1
X_12099_ _01200_ _03482_ _03091_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__or3_1
X_11119_ _04910_ _04907_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__and2_1
Xinput6 data_in[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_2
XFILLER_0_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06660_ _00787_ _00790_ _00732_ VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06591_ result_reg_mac\[2\] VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08330_ _02252_ _02256_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08261_ _02129_ _02189_ _00003_ _02190_ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__a211o_1
X_07212_ _01161_ _01281_ _01294_ VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__a21bo_4
XFILLER_0_74_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08192_ _02123_ _00832_ _02099_ VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_30_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07143_ CMD_set _00697_ _01162_ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__or3_1
XFILLER_0_54_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07074_ _00641_ _00640_ _00654_ _00530_ _01158_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__o311a_4
XFILLER_0_100_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07976_ _01242_ _01247_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__nand2_2
X_06927_ result_reg_not\[13\] VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__inv_2
X_09715_ _03612_ _03616_ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09646_ _03554_ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__inv_2
X_06858_ result_reg_add\[11\] VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06789_ result_reg_set\[8\] _00608_ _00601_ _00915_ VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__o211a_1
X_09577_ _02992_ Qset\[1\]\[6\] _02991_ VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__a21o_1
X_08528_ _02373_ H\[0\]\[12\] VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08459_ _02376_ _02380_ _01553_ VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__a21o_2
XFILLER_0_92_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11470_ _05361_ _05370_ VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__or2_1
X_10421_ _04244_ _04326_ _04239_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__nand3_1
X_10352_ _04257_ _02649_ _02753_ _04258_ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__a211o_1
XFILLER_0_103_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12022_ _05853_ VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__inv_2
X_10283_ _04181_ _04189_ VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12924_ clknet_leaf_17_clk _00367_ VGND VGND VPWR VPWR result_reg_or\[11\] sky130_fd_sc_hd__dfxtp_1
X_12855_ clknet_leaf_18_clk _00298_ VGND VGND VPWR VPWR result_reg_mac\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11806_ result_reg_mul\[6\] _05669_ _05682_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__o21ai_1
X_12786_ clknet_leaf_54_clk _00229_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11737_ _00635_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11668_ _05561_ _05567_ VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11599_ _04835_ _05494_ _05496_ _05498_ VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__o31a_1
X_10619_ _04523_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07830_ result_reg_mul\[13\] _01679_ _01656_ VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__o21ai_1
X_07761_ _00949_ _01608_ _01600_ _01816_ VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__a211o_1
XFILLER_0_47_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06712_ _00841_ _00812_ _00611_ VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__mux2_1
X_09500_ _03408_ _03409_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__nand2_1
X_07692_ result_reg_mul\[6\] _01688_ _01667_ VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06643_ net10 _00600_ _00739_ VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_63_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09431_ _02582_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_35_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06574_ result_reg_or\[1\] VGND VGND VPWR VPWR _00708_ sky130_fd_sc_hd__inv_2
X_09362_ _03267_ _03271_ _03272_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08313_ _02230_ Qset\[2\]\[4\] VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__nand2_1
XANTENNA_22 _00802_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_11 _00677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09293_ _03203_ _03199_ VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__nand2_1
XANTENNA_44 _01085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 _00904_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 _01349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08244_ _02172_ _00003_ _02173_ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__nand3_1
XANTENNA_66 _01437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 _01757_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 _01591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08175_ im_reg\[6\] _02100_ _02105_ _02111_ VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_99 _01819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07126_ _01205_ _01207_ _01208_ _01210_ VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07057_ _01106_ Qset\[2\]\[15\] _01128_ VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07959_ _01964_ VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__inv_2
X_10970_ _04869_ _04870_ _04871_ _04872_ _00621_ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_87_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09629_ _03403_ _03381_ VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12640_ clknet_leaf_54_clk _00090_ VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12571_ clknet_leaf_34_clk _00021_ VGND VGND VPWR VPWR next_PC\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11522_ _05421_ _05422_ VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__nand2_1
X_11453_ _05350_ _05351_ _05352_ _05353_ _00647_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__a221o_1
X_10404_ _04281_ _04309_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__nor2_1
X_11384_ _05109_ _05285_ VGND VGND VPWR VPWR _05286_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10335_ _04240_ _04241_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__or2_1
X_10266_ _03919_ _03921_ _03956_ VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__o21bai_1
X_12005_ _05755_ _05833_ VGND VGND VPWR VPWR _05841_ sky130_fd_sc_hd__nor2_1
X_10197_ _03152_ H\[2\]\[12\] VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_49_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12907_ clknet_leaf_16_clk _00350_ VGND VGND VPWR VPWR result_reg_and\[10\] sky130_fd_sc_hd__dfxtp_1
X_12838_ clknet_leaf_4_clk _00281_ VGND VGND VPWR VPWR result_reg_mul\[5\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_68_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12769_ clknet_leaf_26_clk _00212_ VGND VGND VPWR VPWR H\[0\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_41_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06290_ _06256_ net22 VGND VGND VPWR VPWR _06257_ sky130_fd_sc_hd__nand2_1
Xinput20 instruction_in[12] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_1
XFILLER_0_71_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput31 instruction_in[6] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09980_ _02619_ _03876_ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_52 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08931_ Oset\[1\]\[2\] _02688_ _02840_ VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__a21o_1
X_08862_ _02773_ _02774_ VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__nand2_1
X_07813_ _01863_ _01658_ _01864_ _01865_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__a31o_1
X_08793_ _02705_ _00007_ _02706_ VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__nand3_1
X_07744_ _01797_ _01800_ _01613_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__mux2_2
XFILLER_0_74_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07675_ _01594_ _01727_ _01734_ VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__o21ai_1
X_06626_ _00664_ _00751_ _00758_ VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__o21ai_4
X_09414_ _03323_ VGND VGND VPWR VPWR _03324_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06557_ result_reg_Lshift\[1\] VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09345_ _03254_ _03255_ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_32_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06488_ _00622_ VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__clkbuf_4
X_09276_ _03182_ _03148_ _03149_ VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08227_ _02154_ _02157_ _01551_ VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__a21o_2
X_08158_ _01148_ VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__buf_4
X_07109_ net1 _01193_ VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__nor2_1
X_08089_ _01700_ H\[1\]\[3\] _02057_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10120_ _04024_ _04026_ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__nand2_1
X_10051_ _03942_ _03924_ VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_89_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10953_ _04855_ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10884_ _04786_ _03048_ _04787_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__nand3_1
XFILLER_0_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
X_12623_ clknet_leaf_51_clk _00073_ VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12554_ _01054_ Qset\[3\]\[13\] _06233_ VGND VGND VPWR VPWR _06248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11505_ _05404_ _05402_ VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__nand2b_1
X_12485_ _02116_ _06208_ VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__nor2_1
X_11436_ H\[2\]\[14\] H\[3\]\[14\] _05319_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11367_ _05267_ _05268_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_21_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10318_ _04223_ _04224_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__nand2_1
X_11298_ _05197_ _05199_ VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10249_ _04041_ _04155_ VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07460_ _01528_ VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__clkbuf_1
X_07391_ _01208_ _01014_ VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__nand2_1
X_06411_ shift.left CMD_logic_shift_right VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_14_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
X_06342_ next_PC\[2\] _00481_ VGND VGND VPWR VPWR _00485_ sky130_fd_sc_hd__or2_1
X_09130_ _03022_ Oset\[2\]\[4\] VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__nand2_1
X_09061_ Oset\[3\]\[3\] _02688_ _02837_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__a21oi_1
X_08012_ _02018_ VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__buf_4
XFILLER_0_102_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09963_ _02527_ H\[0\]\[10\] VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__or2_1
X_08914_ _02825_ _02786_ VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__nand2_1
X_09894_ Oset\[0\]\[8\] Oset\[1\]\[8\] _03791_ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__mux2_1
X_08845_ _02585_ Qset\[1\]\[2\] VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__nand2_1
X_08776_ H\[3\]\[1\] _02688_ _02626_ _02689_ VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__a211o_1
X_07727_ result_reg_mul\[8\] _01679_ _01656_ VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07658_ result_reg_not\[4\] _01633_ _01718_ VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_84_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07589_ _00728_ _00729_ _01545_ VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__mux2_1
X_06609_ result_reg_sub\[2\] _00740_ _00741_ VGND VGND VPWR VPWR _00742_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09328_ _02905_ _03238_ VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_51_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09259_ _03169_ _02552_ VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12270_ _06039_ _05812_ _06044_ _06046_ VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11221_ _04636_ VGND VGND VPWR VPWR _05124_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11152_ _04719_ _04716_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__nand2_1
X_10103_ _03987_ _04009_ VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__nand2_1
X_11083_ _04495_ _04975_ _04985_ VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__or3_1
X_10034_ _03924_ _03938_ _03940_ VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_59_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11985_ _05824_ VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10936_ _04838_ _03760_ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__nand2_1
X_10867_ _04764_ _04770_ VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12606_ clknet_leaf_49_clk _00056_ VGND VGND VPWR VPWR Qset\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10798_ _04648_ _04698_ _04701_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_26_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12537_ _06239_ VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__clkbuf_1
X_12468_ _06196_ _06123_ _06267_ VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11419_ _05319_ _02483_ VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__nor2_1
X_12399_ _06116_ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06960_ _01080_ Qset\[0\]\[14\] _00686_ VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_3_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
X_06891_ result_reg_or\[12\] VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__inv_2
X_08630_ _02544_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__buf_4
XFILLER_0_55_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08561_ _02459_ Qset\[3\]\[14\] _02374_ _02477_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07512_ _00557_ _00631_ _00634_ _01576_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__or4_4
XFILLER_0_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08492_ _02408_ _02411_ VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__nand2_2
X_07443_ result_reg_add\[15\] _01267_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07374_ _00991_ _00982_ _01174_ VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09113_ _02836_ VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__buf_2
XFILLER_0_72_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06325_ R3\[0\] _06285_ VGND VGND VPWR VPWR _00470_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_20_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09044_ _02955_ _02828_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09946_ _02372_ _02565_ _03135_ _03852_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__a211o_1
X_09877_ _03782_ _03783_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08828_ _00622_ _02735_ _02741_ VGND VGND VPWR VPWR _02742_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_56_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ _02672_ VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__inv_2
X_11770_ _05132_ _05133_ _05655_ _05656_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__a31o_1
XFILLER_0_67_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10721_ _04622_ _04623_ _03794_ _04624_ _04625_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__a32o_1
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10652_ _04347_ _04556_ VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10583_ _04283_ H\[0\]\[10\] VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12322_ R3\[0\] _05744_ _00498_ _05745_ _06054_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__a221o_1
XFILLER_0_51_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12253_ _06033_ _00778_ VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11204_ _05106_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12184_ _03128_ _03328_ _05892_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11135_ _05036_ _05037_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__or2_1
X_11066_ _04966_ _04968_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10017_ _03923_ VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11968_ _01554_ _03874_ VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11899_ _00589_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__clkbuf_4
X_10919_ _04816_ _04819_ _04633_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__nand3_1
XFILLER_0_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_22 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07090_ _00610_ _00542_ _01174_ VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09800_ _03707_ _00831_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__nand2_1
X_07992_ _02008_ VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__clkbuf_1
X_06943_ _00714_ result_reg_or\[14\] VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__nand2_1
X_09731_ _03635_ _03636_ _03637_ _03638_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__o22a_2
X_06874_ _00981_ _00695_ _00997_ _00725_ _00644_ VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__a221o_1
X_09662_ _03569_ _00623_ _03570_ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__nand3_1
X_09593_ _03345_ _03497_ _03499_ _03501_ VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__a31o_2
X_08613_ _02527_ VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__buf_6
XFILLER_0_89_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08544_ _02459_ Oset\[3\]\[13\] _02374_ _02461_ VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_53_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08475_ H\[3\]\[10\] VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07426_ net6 _01193_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07357_ result_reg_mul\[10\] _01263_ _01245_ _01431_ VGND VGND VPWR VPWR _01432_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_33_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06308_ _06270_ VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07288_ _01358_ _01214_ _01365_ _01159_ _01366_ VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__a311o_1
XFILLER_0_60_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09027_ _02592_ _02231_ VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_79_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_68_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09929_ Qset\[3\]\[9\] _03136_ VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12940_ clknet_leaf_21_clk _00383_ VGND VGND VPWR VPWR result_reg_not\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_5_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ clknet_leaf_23_clk _00314_ VGND VGND VPWR VPWR result_reg_Lshift\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _01830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_134 _06012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11822_ result_reg_mul\[11\] _05670_ _05672_ _05693_ VGND VGND VPWR VPWR _00287_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_123 _04721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 _02168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_167 _00997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_145 im_reg\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_156 R2\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11753_ _05627_ _03740_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_178 _01905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_189 _00809_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10704_ _04606_ _04608_ VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__nand2_1
X_11684_ _05574_ _05583_ VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__xor2_1
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10635_ _03874_ VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12305_ _06058_ _06069_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__nand2_1
X_10566_ _02395_ _02162_ VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_86_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10497_ _04401_ _04196_ _04402_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__nand3_1
X_12236_ _06024_ _01243_ _05338_ _01666_ _05947_ VGND VGND VPWR VPWR _06025_ sky130_fd_sc_hd__a221o_1
X_12167_ result_reg_or\[1\] _05959_ _05967_ _05968_ _05940_ VGND VGND VPWR VPWR _00357_
+ sky130_fd_sc_hd__o221a_1
X_11118_ _05011_ _05020_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__xor2_1
X_12098_ result_reg_and\[5\] _05894_ _05908_ _05911_ _02125_ VGND VGND VPWR VPWR _00345_
+ sky130_fd_sc_hd__o221a_1
Xinput7 data_in[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_2
X_11049_ _04950_ _04897_ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06590_ _00723_ VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08260_ H\[1\]\[1\] _02129_ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__nor2_1
X_07211_ _00724_ _01220_ _01160_ _01293_ VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__a211o_1
X_08191_ _02121_ _02122_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07142_ _01226_ _01214_ VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07073_ _01157_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__buf_4
XFILLER_0_42_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07975_ _01986_ _01998_ _01996_ LC\[9\] VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__a22o_1
X_06926_ _01031_ _00695_ _01047_ _00725_ _00644_ VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__a221o_1
X_09714_ _03504_ _02308_ _03303_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06857_ result_reg_mac\[11\] VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_2_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09645_ _03552_ _03542_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_66_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06788_ _00914_ _00615_ VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__nand2_1
X_09576_ _02992_ _02292_ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08527_ H\[1\]\[12\] VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08458_ _02377_ _02373_ _02378_ _02379_ VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__a211o_1
X_07409_ _01480_ _01255_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10420_ _04324_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__inv_2
X_08389_ _02241_ _02312_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10351_ result_reg_add\[8\] _02648_ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10282_ _04187_ _04188_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12021_ _05770_ _05851_ _05775_ _05852_ VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__a211o_1
X_12923_ clknet_leaf_17_clk _00366_ VGND VGND VPWR VPWR result_reg_or\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12854_ clknet_leaf_18_clk _00297_ VGND VGND VPWR VPWR result_reg_mac\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11805_ _00472_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__clkbuf_4
X_12785_ clknet_leaf_54_clk _00228_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dfxtp_1
X_11736_ _05633_ VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11667_ _05565_ _05566_ VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_94_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11598_ _05335_ Oset\[3\]\[15\] _04303_ _05497_ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__a211o_1
X_10618_ _04520_ _04522_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10549_ _04449_ _04453_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12219_ _03866_ _04671_ _01666_ VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07760_ result_reg_Rshift\[9\] _01608_ VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__nor2_1
X_06711_ result_reg_sub\[5\] VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07691_ _01579_ result_reg_sub\[6\] VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__nand2_1
X_09430_ _03339_ _02556_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__nand2_1
X_06642_ result_reg_set\[3\] _00615_ _00696_ _00773_ VGND VGND VPWR VPWR _00774_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_63_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06573_ net8 _00696_ _00699_ _00706_ VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09361_ _03224_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08312_ _02239_ VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__clkbuf_1
X_09292_ _03148_ _03109_ VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__nand2_1
XANTENNA_23 _00814_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_12 _00677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08243_ _02127_ Qset\[3\]\[1\] VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__nand2_1
XANTENNA_34 _00909_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_45 _01098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_56 _01349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_89 _01768_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08174_ _02102_ _02103_ net44 VGND VGND VPWR VPWR _02111_ sky130_fd_sc_hd__a21o_1
XANTENNA_78 _01621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_67 _01437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07125_ _01209_ _01207_ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__nor2_1
X_07056_ _01144_ VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07958_ _01985_ VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__clkbuf_1
X_06909_ result_reg_mac\[13\] VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__inv_2
X_07889_ _01938_ H\[3\]\[15\] _01628_ VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09628_ _03230_ _03406_ _03231_ VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__nand3_1
X_09559_ _03463_ _03301_ VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__nand2_1
X_12570_ clknet_leaf_36_clk _00020_ VGND VGND VPWR VPWR next_PC\[6\] sky130_fd_sc_hd__dfxtp_1
X_11521_ _05420_ _05414_ VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__nand2_1
X_11452_ Oset\[1\]\[14\] _04858_ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10403_ _04308_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__clkinv_4
X_11383_ _05088_ _05105_ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__or2_1
X_10334_ _03681_ _03674_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10265_ _04169_ _04171_ VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__nand2_1
X_12004_ result_reg_Lshift\[14\] _05743_ _05808_ _05840_ VGND VGND VPWR VPWR _00322_
+ sky130_fd_sc_hd__o211a_1
X_10196_ H\[0\]\[12\] H\[1\]\[12\] _02567_ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12906_ clknet_leaf_17_clk _00349_ VGND VGND VPWR VPWR result_reg_and\[9\] sky130_fd_sc_hd__dfxtp_1
X_12837_ clknet_leaf_56_clk _00280_ VGND VGND VPWR VPWR result_reg_mul\[4\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_83_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12768_ clknet_leaf_33_clk _00211_ VGND VGND VPWR VPWR H\[0\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12699_ clknet_leaf_29_clk _00149_ VGND VGND VPWR VPWR Oset\[0\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_11719_ _05617_ _05618_ VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput10 data_in[3] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
Xinput21 instruction_in[13] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput32 instruction_in[7] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08930_ Oset\[2\]\[2\] Oset\[3\]\[2\] _02688_ VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__mux2_1
X_08861_ _02206_ _00583_ VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__nand2_1
X_07812_ net4 _01746_ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08792_ _02527_ Qset\[3\]\[1\] VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__nand2_1
X_07743_ result_reg_not\[8\] _01633_ _01799_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07674_ _01731_ _01572_ _01732_ _01568_ _01733_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__a311o_1
X_06625_ _00752_ _00655_ _00657_ _00757_ _00666_ VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__a221o_2
X_09413_ _02582_ Qset\[0\]\[5\] VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06556_ result_reg_Rshift\[1\] VGND VGND VPWR VPWR _00690_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09344_ _03252_ _03244_ _03249_ VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__nand3_1
XFILLER_0_62_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06487_ CMD_mul_accumulation VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__clkbuf_4
X_09275_ _03185_ VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08226_ _02151_ _02155_ _02143_ _02156_ VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__a211o_1
XFILLER_0_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08157_ _02095_ _02099_ VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__nand2_4
X_07108_ _01186_ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__buf_2
XFILLER_0_15_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08088_ _02060_ VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07039_ _00878_ Qset\[2\]\[6\] _01129_ VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10050_ _03922_ _03944_ _03956_ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_89_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10952_ _04415_ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10883_ _04600_ _04784_ _04597_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__nand3_1
X_12622_ clknet_leaf_1_clk _00072_ VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__dfxtp_1
X_12553_ _06247_ VGND VGND VPWR VPWR _00464_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11504_ _05402_ _05404_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_80_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12484_ _06102_ _00620_ _06117_ _06124_ VGND VGND VPWR VPWR _06208_ sky130_fd_sc_hd__o22a_1
X_11435_ _02494_ _05335_ _04835_ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11366_ _05266_ _05258_ VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__nand2_1
X_10317_ _03662_ _03659_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__or2_1
X_11297_ _05198_ _05027_ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__nand2_1
X_10248_ _04152_ _04154_ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_13_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10179_ _04082_ _04083_ _04084_ _04085_ VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__a22o_2
XFILLER_0_88_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06410_ CMD_or VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07390_ _01459_ _01462_ _01271_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06341_ _00481_ next_PC\[2\] VGND VGND VPWR VPWR _00484_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09060_ _02968_ _02969_ _02970_ _02971_ Oreg3 VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__a221o_1
X_08011_ _01225_ _01999_ VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__nor2_4
XFILLER_0_25_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09962_ _02785_ _03868_ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_31_Left_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08913_ _02786_ _02825_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__or2_1
X_09893_ H\[1\]\[8\] _03793_ _03798_ _03799_ VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__a211o_1
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08844_ _02581_ Qset\[0\]\[2\] VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__nand2_1
X_08775_ _02688_ _02186_ VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__nor2_1
X_07726_ _00912_ _00906_ _01545_ VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07657_ result_reg_Rshift\[4\] _01672_ _01607_ _01717_ VGND VGND VPWR VPWR _01718_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06608_ _00540_ _00729_ _00534_ VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__a21oi_1
X_07588_ _01651_ VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06539_ _00672_ _00628_ _00664_ _00673_ VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__a211o_1
X_09327_ _02785_ _02821_ VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_51_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09258_ _02560_ _03164_ _03166_ _03168_ VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_50_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09189_ _02874_ H\[3\]\[6\] _02534_ VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08209_ _02139_ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__buf_8
X_11220_ _04820_ _04633_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_95_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11151_ _04953_ _04196_ _05053_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__nand3_1
X_10102_ _04008_ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__inv_2
X_11082_ _04958_ _04983_ _04984_ VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__o21ai_1
X_10033_ _03939_ _03925_ VGND VGND VPWR VPWR _03940_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11984_ _05822_ _05771_ _05775_ _05823_ VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__a211o_1
XFILLER_0_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10935_ Oset\[3\]\[12\] VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10866_ _04765_ _04769_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_104_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12605_ clknet_leaf_25_clk _00055_ VGND VGND VPWR VPWR Qset\[1\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_10797_ _04507_ _04700_ VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12536_ _00809_ Qset\[3\]\[4\] _06234_ VGND VGND VPWR VPWR _06239_ sky130_fd_sc_hd__mux2_1
X_12467_ _06178_ _06157_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11418_ _04832_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__buf_2
XFILLER_0_34_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12398_ _06138_ VGND VGND VPWR VPWR _06139_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11349_ _05087_ _05083_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06890_ _01009_ _00743_ _01011_ _01012_ VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__a31o_1
X_13019_ clknet_leaf_35_clk _00462_ VGND VGND VPWR VPWR Qset\[3\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_08560_ _02459_ _02476_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__nor2_1
X_07511_ shift.left CMD_logic_shift_right _00624_ _01575_ VGND VGND VPWR VPWR _01576_
+ sky130_fd_sc_hd__or4_1
XFILLER_0_49_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08491_ _02328_ Qset\[1\]\[11\] _02329_ _02410_ VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__a211o_1
X_07442_ result_reg_and\[15\] _01299_ VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07373_ result_reg_set\[11\] VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__inv_2
X_06324_ _06284_ VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__buf_2
X_09112_ _03022_ VGND VGND VPWR VPWR _03023_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09043_ _02951_ _02953_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09945_ _02565_ H\[2\]\[9\] VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__nor2_1
X_09876_ _02341_ _02162_ VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__nand2_1
X_08827_ _02737_ _00622_ _02740_ VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_56_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _02671_ _01153_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__nand2_1
X_07709_ result_reg_mul\[7\] _01653_ _01561_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08689_ _02602_ _02590_ _02603_ VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__nand3_4
X_10720_ _03023_ Oset\[2\]\[10\] VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10651_ _03790_ _04555_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__nand2_1
X_10582_ H\[2\]\[10\] H\[3\]\[10\] _04282_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12321_ _06079_ _06080_ _02125_ VGND VGND VPWR VPWR _00399_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12252_ _06032_ _05753_ _06013_ _06036_ VGND VGND VPWR VPWR _00374_ sky130_fd_sc_hd__o211a_1
X_11203_ _05088_ _05105_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__xnor2_1
X_12183_ result_reg_or\[4\] _05959_ _05857_ _05981_ VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11134_ _04309_ _04899_ _05020_ _05018_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__o31a_1
X_11065_ _04881_ Oset\[3\]\[13\] _04045_ _04967_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__a211o_1
X_10016_ _03902_ _03895_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__nand2_1
X_11967_ _05774_ _05807_ _05808_ _05809_ VGND VGND VPWR VPWR _00316_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10918_ _04820_ _04821_ VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11898_ _05744_ _02538_ _05745_ _02550_ _05747_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__a221o_2
X_10849_ _04751_ _04752_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12519_ next_PC\[7\] _06218_ VGND VGND VPWR VPWR _06229_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07991_ Oset\[0\]\[6\] _01368_ _02001_ VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_105_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06942_ _01059_ _00562_ _01061_ _01062_ VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__a31o_1
XFILLER_0_66_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09730_ Qset\[1\]\[7\] _03341_ _03004_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__o21ai_1
X_06873_ _00739_ _00988_ _00990_ _00995_ _00996_ VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__a32o_1
X_09661_ _03562_ _03563_ _03233_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__nand3_1
X_08612_ _00006_ VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__buf_6
X_09592_ _02992_ _02303_ _03004_ _03500_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__o211a_1
X_08543_ _02459_ _02460_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_81_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08474_ _02392_ _02393_ _02394_ _02378_ VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__a22oi_4
X_07425_ _01066_ _01495_ _01181_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07356_ result_reg_add\[10\] _01264_ _01266_ _01430_ VGND VGND VPWR VPWR _01431_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_33_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07287_ result_reg_mac\[6\] _01215_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__nor2_1
X_06307_ _06269_ _06261_ VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09026_ _02936_ _02937_ VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_79_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09928_ _03833_ _03834_ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_69_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09859_ _03760_ H\[1\]\[8\] _03764_ _03765_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__a211o_1
X_12870_ clknet_leaf_23_clk _00313_ VGND VGND VPWR VPWR result_reg_Lshift\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_102 _01834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_124 _05115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11821_ _04722_ _04791_ _05673_ VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__a21o_1
XANTENNA_113 _02382_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_135 _06030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_146 im_reg\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_157 R2\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11752_ _05644_ VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_168 _01047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_179 _02101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _04607_ _02096_ VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__nand2_1
X_11683_ _05581_ _05582_ _04196_ VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__a21oi_1
X_10634_ _04345_ _04309_ VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12304_ _00681_ _02311_ _03094_ _02139_ _03105_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__o221a_1
X_10565_ _04463_ _04469_ _04464_ VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__nand3_1
X_10496_ _04364_ _04366_ _03048_ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__a21o_1
X_12235_ _05324_ _04064_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__nand2_1
X_12166_ _05904_ _02682_ _05884_ _05957_ VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__a211o_1
X_11117_ _05018_ _05019_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__nand2_1
X_12097_ _05888_ _03141_ _03346_ _05910_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__o31ai_1
Xinput8 data_in[1] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dlymetal6s2s_1
X_11048_ _04897_ _04950_ VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12999_ clknet_leaf_39_clk _00442_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07210_ _01287_ _01292_ _01214_ VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__and3_1
X_08190_ _00597_ CMD_store _00697_ VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__nand3_1
XFILLER_0_15_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07141_ R1\[1\] VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07072_ _00589_ _01156_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__nor2_2
XFILLER_0_2_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07974_ _01997_ im_reg\[9\] _01960_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06925_ _01040_ _00619_ _01046_ VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__a21o_1
X_09713_ _03620_ _03459_ VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09644_ _03542_ _03552_ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__nor2_1
X_06856_ _00980_ VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_66_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06787_ _00911_ _00913_ _00613_ VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__mux2_1
X_09575_ _03483_ VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08526_ _02443_ _02444_ VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08457_ _02373_ H\[0\]\[9\] VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__nor2_1
X_07408_ _01033_ _01479_ _01182_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08388_ Qset\[2\]\[7\] VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07339_ _00930_ _01414_ _01181_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__mux2_1
X_10350_ _04256_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10281_ _04010_ _04182_ _04185_ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__nand3_1
X_09009_ _02585_ Oset\[1\]\[3\] VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12020_ result_reg_Rshift\[3\] _05851_ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__nor2_1
X_12922_ clknet_leaf_17_clk _00365_ VGND VGND VPWR VPWR result_reg_or\[9\] sky130_fd_sc_hd__dfxtp_1
X_12853_ clknet_leaf_18_clk _00296_ VGND VGND VPWR VPWR result_reg_mac\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12784_ clknet_leaf_2_clk _00227_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dfxtp_1
X_11804_ _05681_ VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11735_ _00702_ _05628_ _02753_ _05632_ VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__a211o_1
XFILLER_0_83_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11666_ _05564_ _03145_ _04494_ _04196_ VGND VGND VPWR VPWR _05566_ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11597_ _05335_ _02507_ VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__nor2_1
X_10617_ _04516_ _04521_ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__nand2_1
X_10548_ _04450_ _04451_ _04452_ VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_24_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12218_ _04741_ _04677_ _05892_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__a21oi_1
X_10479_ _04383_ _04384_ VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__nand2_1
X_12149_ _05515_ _05951_ _05499_ _05952_ VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06710_ result_reg_set\[5\] VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__inv_2
X_07690_ _01580_ result_reg_add\[6\] VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__nand2_1
X_06641_ _00772_ _00615_ VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06572_ _00700_ _00705_ _00607_ VGND VGND VPWR VPWR _00706_ sky130_fd_sc_hd__mux2_1
X_09360_ _03269_ _03270_ VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__nand2_1
X_08311_ _02238_ net57 _02170_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__mux2_1
X_09291_ _03200_ _03201_ VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__nand2_1
XANTENNA_13 _00683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08242_ _02128_ Qset\[2\]\[1\] VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__nand2_1
XANTENNA_57 _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 _00946_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 _00818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 _01149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_79 _01668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_68 _01444_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08173_ R1\[1\] _02100_ _02105_ _02110_ VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__o211a_1
X_07124_ result_reg_and\[0\] VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07055_ _01080_ Qset\[2\]\[14\] _01128_ VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07957_ _01984_ LC\[5\] _01964_ VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__mux2_1
X_06908_ _01030_ VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07888_ _01934_ _01937_ _01612_ VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06839_ net2 _00696_ _00963_ VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__o21ai_1
X_09627_ _03535_ _03274_ VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_87_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09558_ _03459_ _03464_ VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__nand2_1
X_08509_ _02428_ VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11520_ _05414_ _05420_ VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__or2_1
X_09489_ _03397_ _03398_ VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11451_ _04855_ Oset\[0\]\[14\] _04862_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__a21oi_1
X_11382_ _05283_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__inv_2
X_10402_ _04307_ _02381_ VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__nand2_8
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10333_ _04237_ _04239_ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10264_ _04112_ _04147_ _04170_ VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__o21ai_1
X_12003_ _05839_ _05771_ VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__nand2_1
X_10195_ _04100_ _04101_ VGND VGND VPWR VPWR _04102_ sky130_fd_sc_hd__nand2_1
X_12905_ clknet_leaf_31_clk _00348_ VGND VGND VPWR VPWR result_reg_and\[8\] sky130_fd_sc_hd__dfxtp_2
X_12836_ clknet_leaf_7_clk _00279_ VGND VGND VPWR VPWR result_reg_mul\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12767_ clknet_leaf_33_clk _00210_ VGND VGND VPWR VPWR H\[0\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_11718_ _05613_ _05614_ _05476_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__nand3_1
X_12698_ clknet_leaf_34_clk _00148_ VGND VGND VPWR VPWR Oset\[0\]\[12\] sky130_fd_sc_hd__dfxtp_1
Xinput11 data_in[4] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
Xinput22 instruction_in[14] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
XFILLER_0_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11649_ _05548_ _05048_ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput33 instruction_in[8] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08860_ _02763_ _02772_ VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__nand2_1
X_07811_ _01465_ _01682_ VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__or2_1
X_08791_ _02522_ Qset\[2\]\[1\] VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__nand2_1
X_07742_ result_reg_Rshift\[8\] _01672_ _01607_ _01798_ VGND VGND VPWR VPWR _01799_
+ sky130_fd_sc_hd__o211a_1
X_07673_ result_reg_or\[5\] _01595_ VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_48_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06624_ result_reg_Rshift\[2\] _00753_ _00756_ VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09412_ _03321_ _02591_ VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__nand2_1
X_09343_ _03250_ _03253_ VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__nand2_1
X_06555_ result_reg_not\[1\] VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__inv_2
X_06486_ Oreg3 VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_7_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09274_ _03176_ _03184_ VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08225_ H\[1\]\[0\] _02151_ VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__nor2_1
X_08156_ _00557_ _02098_ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__nor2_4
X_07107_ _01191_ VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08087_ _01676_ H\[1\]\[2\] _02057_ VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07038_ _01135_ VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_89_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08989_ _02785_ _02734_ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10951_ _04853_ _02449_ VGND VGND VPWR VPWR _04854_ sky130_fd_sc_hd__nand2_8
X_12621_ clknet_leaf_27_clk _00071_ VGND VGND VPWR VPWR Qset\[2\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_10882_ _04723_ _04785_ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__nand2_1
X_12552_ _01029_ Qset\[3\]\[12\] _06233_ VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12483_ _06102_ Qreg2 _06206_ _06207_ _02101_ VGND VGND VPWR VPWR _00434_ sky130_fd_sc_hd__o221a_1
X_11503_ _04178_ _05403_ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11434_ _05319_ VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__buf_2
XFILLER_0_61_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11365_ _05258_ _05266_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10316_ _03666_ _03606_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__nand2_1
X_11296_ _05026_ _05010_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__or2_1
X_10247_ _04138_ _04153_ _04139_ VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__nand3b_1
X_10178_ _02545_ Oset\[1\]\[15\] VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_17_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12819_ clknet_leaf_11_clk _00262_ VGND VGND VPWR VPWR result_reg_sub\[2\] sky130_fd_sc_hd__dfxtp_1
X_06340_ _00479_ _00475_ _00483_ next_PC\[1\] _00478_ VGND VGND VPWR VPWR _00015_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_29_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08010_ _02017_ VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09961_ _03867_ VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__buf_4
X_08912_ _02739_ _02822_ _02824_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09892_ _03792_ _02350_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08843_ _02754_ _02584_ _02755_ VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__nand3_1
X_08774_ _02625_ VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07725_ _01782_ VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__clkbuf_1
X_07656_ _01716_ _00806_ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_84_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06607_ _00540_ VGND VGND VPWR VPWR _00740_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07587_ _01650_ H\[3\]\[1\] _01629_ VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__mux2_1
X_06538_ R1\[1\] _00628_ VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__nor2_1
X_09326_ _03235_ _02950_ _03236_ VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09257_ _03157_ Oset\[3\]\[4\] _02535_ _03167_ VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__a211o_1
XFILLER_0_105_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06469_ result_reg_or\[0\] _00553_ result_reg_and\[0\] _00562_ _00603_ VGND VGND
+ VPWR VPWR _00604_ sky130_fd_sc_hd__o221a_1
X_08208_ _01162_ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__buf_8
X_09188_ _02562_ H\[1\]\[6\] VGND VGND VPWR VPWR _03099_ sky130_fd_sc_hd__nand2_1
X_08139_ H\[0\]\[11\] _01859_ _02074_ VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11150_ _05051_ _05052_ _03048_ VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__a21o_1
X_10101_ _04006_ _04007_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__nand2_1
X_11081_ _04308_ _04957_ _03790_ _04982_ VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__a22o_1
X_10032_ _03937_ _03935_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_59_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11983_ result_reg_Lshift\[11\] _05741_ VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__nor2_1
X_10934_ _03773_ _02436_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__nand2_1
X_10865_ _04767_ _04768_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_104_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12604_ clknet_leaf_25_clk _00054_ VGND VGND VPWR VPWR Qset\[1\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10796_ _04699_ _04697_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__nor2_1
X_12535_ _06238_ VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12466_ _06191_ _06167_ _06106_ VGND VGND VPWR VPWR _06195_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11417_ _05318_ VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__inv_2
X_12397_ net24 _06253_ VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__nor2_1
X_11348_ _05248_ _05249_ VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__and2_1
X_11279_ _05179_ _05180_ VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__and2b_1
X_13018_ clknet_leaf_39_clk _00461_ VGND VGND VPWR VPWR Qset\[3\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07510_ _01571_ CMD_and VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__nand2_1
X_08490_ _02319_ _02409_ VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__nor2_1
X_07441_ result_reg_not\[15\] _01510_ _01167_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__mux2_1
X_07372_ _01208_ _00989_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06323_ LC\[9\] _06283_ CMD_loopjump VGND VGND VPWR VPWR _06284_ sky130_fd_sc_hd__o21ai_4
X_09111_ _03021_ VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09042_ _02863_ _02951_ _02953_ VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__nand3_1
XFILLER_0_4_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09944_ H\[1\]\[9\] _03152_ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__nor2_1
X_09875_ _03780_ _00582_ _03781_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__a21oi_1
X_08826_ _02578_ _02738_ _02739_ VGND VGND VPWR VPWR _02740_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_56_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08757_ _02667_ _02670_ _02551_ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__nand3_1
X_07708_ _00883_ _00884_ _01545_ VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08688_ _02585_ Oset\[1\]\[0\] VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07639_ _01700_ H\[3\]\[3\] _01629_ VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__mux2_1
X_10650_ _03768_ _04540_ _04554_ _02811_ _00589_ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09309_ _03145_ _03080_ VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10581_ _02390_ _00585_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12320_ _05766_ _06061_ VGND VGND VPWR VPWR _06080_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12251_ _06033_ _00752_ VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__nand2_1
X_11202_ _05103_ _05104_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12182_ _05937_ _05978_ _05979_ _05980_ _05957_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_101_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11133_ _05029_ _05035_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__xor2_1
X_11064_ _04881_ _02460_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__nor2_1
X_10015_ _03919_ _03921_ VGND VGND VPWR VPWR _03922_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11966_ _05774_ _00923_ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__nand2_1
X_10917_ _04633_ VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__inv_2
X_11897_ _01554_ _05746_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__nor2_1
X_10848_ _04750_ _04726_ VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10779_ _04679_ _04680_ _04681_ _04682_ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__o22a_2
XFILLER_0_26_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12518_ net71 _06220_ _06221_ _06228_ VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__o211a_1
X_12449_ _06132_ _06112_ VGND VGND VPWR VPWR _06181_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07990_ _02007_ VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06941_ result_reg_and\[14\] _00562_ _00709_ VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09660_ _03529_ _03534_ _03274_ VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__nand3_1
X_06872_ net3 _00600_ _00739_ VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__a21oi_1
X_08611_ _02525_ VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09591_ _03001_ H\[1\]\[6\] VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08542_ Oset\[2\]\[13\] VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_53_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08473_ Qset\[2\]\[10\] Qset\[3\]\[10\] _02319_ VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__mux2_1
X_07424_ _01060_ _01494_ _01176_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07355_ _01264_ _00958_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_61_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07286_ _01363_ _01271_ _01190_ _01364_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__a211o_1
X_06306_ current_state\[6\] VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09025_ _02229_ _00583_ _02571_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_92_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09927_ _00588_ im_reg\[8\] VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_5_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09858_ _03760_ _02350_ VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_69_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _03695_ _03696_ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__nand2_1
X_08809_ _02722_ VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__inv_2
XANTENNA_103 _01850_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_125 _05115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11820_ _05692_ VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__inv_2
XANTENNA_114 _02427_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11751_ _00865_ _05631_ _05634_ _05643_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_147 result_reg_mac\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_136 _06182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_158 R2\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_169 _01285_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10702_ _04555_ VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_101_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11682_ _05580_ _05577_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10633_ _04349_ _04348_ _04353_ VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__o21a_1
X_10564_ _04467_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__inv_2
X_12303_ result_reg_set\[5\] _06063_ _06066_ _06068_ VGND VGND VPWR VPWR _00393_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10495_ _04399_ _03048_ _04400_ VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__nand3_1
X_12234_ _05958_ _06022_ VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__nand2_1
X_12165_ _00524_ _05965_ _05966_ _05937_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__a22o_1
X_11116_ _05017_ _05016_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__nand2_1
X_12096_ _05881_ _03122_ _05909_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__or3b_1
X_11047_ _04949_ VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__inv_2
Xinput9 data_in[2] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_86_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12998_ clknet_leaf_54_clk _00441_ VGND VGND VPWR VPWR R3\[0\] sky130_fd_sc_hd__dfxtp_4
X_11949_ _05779_ _05793_ _05755_ VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07140_ R3\[0\] _01219_ _01224_ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_30_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07071_ _01155_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07973_ LC\[9\] _06283_ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__nor2_1
X_09712_ _03348_ _02286_ _03613_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__a21oi_1
X_06924_ _01041_ _00709_ _00714_ _01045_ _00603_ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_2_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09643_ _03543_ _03551_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__xor2_1
X_06855_ _00979_ Qset\[0\]\[10\] _00686_ VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09574_ _02540_ _03482_ _01154_ VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__o21ai_1
X_06786_ _00912_ _00906_ _00611_ VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__mux2_1
X_08525_ _02378_ VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08456_ _02329_ VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__buf_4
XFILLER_0_37_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07407_ _01034_ _01478_ _01177_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__mux2_1
X_08387_ _00591_ VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__buf_8
XFILLER_0_18_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07338_ _00931_ _01413_ _01176_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07269_ _01161_ _01335_ _01348_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__a21bo_4
XFILLER_0_5_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10280_ _04183_ _04186_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09008_ _02581_ Oset\[0\]\[3\] VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12921_ clknet_leaf_31_clk _00364_ VGND VGND VPWR VPWR result_reg_or\[8\] sky130_fd_sc_hd__dfxtp_2
X_12852_ clknet_leaf_18_clk _00295_ VGND VGND VPWR VPWR result_reg_mac\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12783_ clknet_leaf_28_clk _00226_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dfxtp_4
X_11803_ _03416_ _03417_ _05670_ _05680_ VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_53_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11734_ _05631_ _02750_ VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11665_ _03145_ _04494_ _05564_ VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__a21oi_1
X_10616_ _04519_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11596_ _05495_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10547_ _04318_ _04321_ _04319_ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__nand3_1
X_10478_ _04132_ _04134_ _04131_ VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__a21oi_1
X_12217_ _04735_ _04683_ VGND VGND VPWR VPWR _06009_ sky130_fd_sc_hd__nand2_1
X_12148_ _05881_ _04086_ VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__nor2_1
X_12079_ _05881_ _02923_ _02881_ VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06640_ _00765_ _00771_ _00732_ VGND VGND VPWR VPWR _00772_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06571_ _00701_ _00704_ _00613_ VGND VGND VPWR VPWR _00705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_44_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08310_ _02126_ _02222_ _02140_ _02229_ _02237_ VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__o221ai_4
X_09290_ _03146_ _03114_ _03109_ VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__o21a_1
XANTENNA_14 _00717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08241_ _02171_ VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_25 _00820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 _00953_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_47 _01149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_69 _01462_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08172_ _02102_ _02103_ net43 VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__a21o_1
XANTENNA_58 _01368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07123_ _01199_ VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07054_ _01143_ VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07956_ _01962_ _01226_ _01983_ VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__o21ai_1
X_06907_ _01029_ Qset\[0\]\[12\] _00686_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__mux2_1
X_07887_ result_reg_not\[15\] _01600_ _01936_ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__a21o_1
X_06838_ _00962_ _00735_ VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__nand2_1
X_09626_ _03529_ _03534_ VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__nand2_1
X_06769_ _00889_ _00619_ _00629_ _00896_ VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_87_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09557_ _03460_ _03461_ _03465_ VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__nand3_1
X_08508_ _02427_ net50 _02169_ VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__mux2_1
X_09488_ _03392_ _03395_ _03393_ VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_35_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08439_ _02328_ _02360_ VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11450_ _04855_ Oset\[2\]\[14\] VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__nand2_1
X_11381_ _05280_ _05282_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__nand2_1
X_10401_ _04298_ _04299_ _03758_ _04306_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__a31o_2
XFILLER_0_61_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10332_ _04233_ _04238_ _04234_ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__nand3_2
XFILLER_0_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12002_ _05828_ _05838_ _05754_ VGND VGND VPWR VPWR _05839_ sky130_fd_sc_hd__mux2_1
X_10263_ _02738_ _04110_ _04114_ VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__o21ai_1
X_10194_ _04099_ _04052_ VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12904_ clknet_leaf_16_clk _00347_ VGND VGND VPWR VPWR result_reg_and\[7\] sky130_fd_sc_hd__dfxtp_1
X_12835_ clknet_leaf_8_clk _00278_ VGND VGND VPWR VPWR result_reg_mul\[2\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_26_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12766_ clknet_leaf_40_clk _00209_ VGND VGND VPWR VPWR H\[0\]\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_71_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11717_ _05615_ _05616_ VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__nand2_1
X_12697_ clknet_leaf_38_clk _00147_ VGND VGND VPWR VPWR Oset\[0\]\[11\] sky130_fd_sc_hd__dfxtp_1
Xinput12 data_in[5] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_52_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11648_ _05047_ _05043_ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_12_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput23 instruction_in[15] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_2
X_11579_ _05476_ _05479_ VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__nand2_1
Xinput34 instruction_in[9] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07810_ _01861_ _01653_ _01862_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__a21o_1
X_08790_ _00622_ _02687_ _02703_ VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__o21ai_1
X_07741_ _01716_ _00923_ VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07672_ _01691_ result_reg_and\[5\] VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06623_ _00754_ _00755_ VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__nand2_1
X_09411_ _02611_ Qset\[1\]\[5\] VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_17_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
X_09342_ _03252_ VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__inv_2
X_06554_ _00688_ VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06485_ Qreg3 VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09273_ _03051_ _02949_ VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__nor2_1
X_08224_ H\[0\]\[0\] VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__inv_2
X_08155_ _02097_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__inv_2
X_07106_ _01190_ VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08086_ _02059_ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__clkbuf_1
X_07037_ _00854_ Qset\[2\]\[5\] _01129_ VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08988_ _02898_ _02899_ VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__nand2_1
X_07939_ _06273_ LC\[2\] VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__nand2_1
X_10950_ _04852_ _01553_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__nand2_2
X_09609_ _03516_ _03517_ VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__nand2_1
X_10881_ _04784_ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__inv_2
X_12620_ clknet_leaf_27_clk _00070_ VGND VGND VPWR VPWR Qset\[2\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12551_ _06246_ VGND VGND VPWR VPWR _00463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12482_ _06123_ _06189_ _06267_ _06143_ VGND VGND VPWR VPWR _06207_ sky130_fd_sc_hd__a211o_1
X_11502_ _04163_ _04180_ VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__or2b_1
X_11433_ _05319_ H\[0\]\[14\] VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11364_ _05264_ _05265_ VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__nand2_1
X_11295_ _05195_ _05196_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__nand2_1
X_10315_ _04199_ _04221_ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__xor2_1
X_10246_ _04151_ VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10177_ _02523_ Oset\[0\]\[15\] _02525_ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12818_ clknet_leaf_10_clk _00261_ VGND VGND VPWR VPWR result_reg_sub\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12749_ clknet_leaf_40_clk _00192_ VGND VGND VPWR VPWR H\[1\]\[8\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_69_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_6_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
X_09960_ _03866_ _01552_ _02572_ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__and3_1
X_08911_ _02736_ _02823_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__nand2_1
X_09891_ _02840_ VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_75 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08842_ _02592_ Qset\[3\]\[2\] VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__nand2_1
X_08773_ _02686_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__buf_4
XFILLER_0_79_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07724_ _01781_ H\[3\]\[7\] _01629_ VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__mux2_1
X_07655_ _01603_ VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__clkbuf_4
X_06606_ _00603_ VGND VGND VPWR VPWR _00739_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_84_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07586_ _01613_ _01632_ _01634_ _01648_ _01649_ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__a32o_4
XFILLER_0_75_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06537_ _00670_ _00671_ _00602_ VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09325_ _02912_ _02910_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__nor2_1
X_06468_ _00602_ VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09256_ _02545_ _02249_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08207_ _02133_ _02137_ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06399_ _00527_ _00533_ VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__nor2_4
X_09187_ _02787_ H\[0\]\[6\] VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__nand2_1
X_08138_ _02086_ VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08069_ _02049_ VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11080_ _04308_ _04982_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__nand2_1
X_10100_ _04004_ _04001_ _04002_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__nand3_2
XFILLER_0_11_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10031_ _03925_ _03935_ _03937_ VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ _05755_ _05812_ _05765_ _05821_ VGND VGND VPWR VPWR _05822_ sky130_fd_sc_hd__o22a_1
XFILLER_0_105_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10933_ _04831_ _04833_ _04834_ _04835_ VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__a22o_1
X_10864_ _04578_ _04766_ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12603_ clknet_leaf_28_clk _00053_ VGND VGND VPWR VPWR Qset\[1\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_10795_ _04502_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12534_ _00783_ Qset\[3\]\[3\] _06234_ VGND VGND VPWR VPWR _06238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12465_ _06097_ _00585_ _06185_ _06194_ _02101_ VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11416_ _05315_ _02649_ _05316_ _05317_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__a31o_1
X_12396_ _06126_ _06136_ _04827_ _06137_ VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11347_ _05246_ _05245_ VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11278_ _05178_ _04929_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__nand2_1
X_13017_ clknet_leaf_39_clk _00460_ VGND VGND VPWR VPWR Qset\[3\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_10229_ _04131_ _04134_ _04132_ VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_55_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07440_ result_reg_Lshift\[15\] result_reg_Rshift\[15\] _01164_ VGND VGND VPWR VPWR
+ _01510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07371_ _01441_ _01444_ _01271_ VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06322_ _06281_ _06282_ VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__nand2_2
X_09110_ _02632_ VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__buf_2
XFILLER_0_29_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09041_ _02914_ _02915_ _02952_ VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__nand3_1
XFILLER_0_13_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09943_ _02567_ H\[0\]\[9\] VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09874_ _02552_ VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__clkbuf_4
X_08825_ _02620_ _02734_ VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_56_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08756_ _02668_ _02590_ _02669_ VGND VGND VPWR VPWR _02670_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_28_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07707_ _00899_ _01607_ _01764_ VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08687_ _02581_ Oset\[0\]\[0\] VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__nand2_1
X_07638_ _01696_ _01699_ _01613_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__mux2_4
X_07569_ _01600_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09308_ _03187_ _03183_ _03186_ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__nand3_1
XFILLER_0_90_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10580_ _04471_ _03770_ _04478_ _04484_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09239_ _03148_ _03149_ VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__nand2_1
X_12250_ _06032_ _05759_ _06013_ _06035_ VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12181_ _03155_ _03015_ _05888_ VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__a21oi_1
X_11201_ _04696_ _04695_ _04703_ _04704_ VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_101_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11132_ _05033_ _05034_ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11063_ _04881_ Oset\[1\]\[13\] _04042_ _04965_ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__a211o_1
X_10014_ _03920_ VGND VGND VPWR VPWR _03921_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11965_ _01148_ VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10916_ _04816_ _04819_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__nand2_1
X_11896_ _02570_ VGND VGND VPWR VPWR _05746_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10847_ _04726_ _04750_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10778_ Oset\[1\]\[11\] _03341_ _03004_ VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12517_ _06219_ _00506_ VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12448_ _06097_ _05904_ _06179_ _06180_ _02101_ VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__o221a_1
XFILLER_0_41_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12379_ net24 VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__inv_2
X_06940_ _01060_ _00745_ VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__or2_1
X_06871_ result_reg_set\[11\] _00615_ _00696_ _00994_ VGND VGND VPWR VPWR _00995_
+ sky130_fd_sc_hd__o211ai_1
X_08610_ _00007_ VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_19_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09590_ _03498_ H\[3\]\[6\] VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08541_ _02373_ VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__buf_4
XFILLER_0_49_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08472_ Qset\[1\]\[10\] _02327_ _02347_ VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_81_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07423_ _01067_ _01057_ _01173_ VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07354_ result_reg_and\[10\] _01207_ _01261_ VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_61_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07285_ result_reg_or\[6\] _01199_ VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06305_ _06268_ VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_28_Left_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09024_ _02925_ _02935_ VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_92_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09926_ _03827_ _03832_ VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_37_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ _03345_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_69_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ _01153_ _00669_ _02555_ VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__o21ai_1
X_09788_ _03694_ _03693_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__nand2_1
X_08739_ _02647_ VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_104 _01863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_115 _02450_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11750_ _05627_ _03601_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_148 net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_126 _05298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_137 _06218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_159 R2\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10701_ _04527_ _04605_ _00710_ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__nand3_1
XFILLER_0_76_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11681_ _05577_ _05580_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10632_ _04536_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10563_ _04465_ _04467_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12302_ _06063_ _06067_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10494_ _04194_ _04157_ _04397_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__nand3_1
X_12233_ _05329_ _04058_ _05892_ VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__a21o_1
X_12164_ _02719_ _05882_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_55_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12095_ _03333_ _03335_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__and2_1
X_11115_ _05016_ _05017_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__or2_1
X_11046_ _04947_ _04948_ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12997_ clknet_3_0__leaf_clk _00440_ VGND VGND VPWR VPWR R2\[0\] sky130_fd_sc_hd__dfxtp_4
X_11948_ _05792_ VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11879_ result_reg_mac\[13\] _05702_ _05682_ VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_64_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07070_ _01154_ VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__buf_4
XFILLER_0_42_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07972_ _01995_ _01996_ _06282_ _01993_ VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__o22ai_1
X_09711_ _03615_ _03617_ _03618_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__nand3_1
X_06923_ _01042_ _01044_ _00561_ VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__mux2_1
X_06854_ _00664_ _00973_ _00978_ VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_93_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09642_ _03549_ _03550_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__nand2_1
X_06785_ result_reg_sub\[8\] VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09573_ _03478_ _03479_ _03481_ VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_38_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08524_ H\[2\]\[12\] H\[3\]\[12\] _02397_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08455_ H\[1\]\[9\] VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__inv_2
X_07406_ _01035_ _01036_ _01174_ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__mux2_1
X_08386_ _02310_ VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07337_ _00932_ _00933_ _01173_ VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07268_ _01340_ _01214_ _01346_ _01159_ _01347_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__a311o_1
XFILLER_0_5_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07199_ result_reg_and\[2\] VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__inv_2
X_09007_ _02917_ _02584_ _02918_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__nand3_1
X_09909_ _02545_ Qset\[2\]\[8\] _02526_ VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__o21ai_1
X_12920_ clknet_leaf_16_clk _00363_ VGND VGND VPWR VPWR result_reg_or\[7\] sky130_fd_sc_hd__dfxtp_1
X_12851_ clknet_leaf_18_clk _00294_ VGND VGND VPWR VPWR result_reg_mac\[2\] sky130_fd_sc_hd__dfxtp_1
X_11802_ result_reg_mul\[5\] _05677_ _05134_ VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__o21ai_1
X_12782_ clknet_leaf_27_clk _00225_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dfxtp_1
X_11733_ _05627_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__clkbuf_4
X_11664_ _05562_ _05563_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__xor2_1
X_10615_ _04517_ _04519_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__nand2_1
X_11595_ _05335_ Oset\[1\]\[15\] VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10546_ _04239_ VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10477_ _04381_ _04382_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__nand2_1
X_12216_ result_reg_or\[10\] _05960_ _06006_ _06008_ _02101_ VGND VGND VPWR VPWR _00366_
+ sky130_fd_sc_hd__o221a_1
X_12147_ _05888_ _04093_ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__nor2_1
X_12078_ _05878_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11029_ _04928_ _04931_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__or2_1
X_06570_ _00702_ _00703_ _00611_ VGND VGND VPWR VPWR _00704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08240_ _02159_ net48 _02170_ VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__mux2_1
XANTENNA_26 _00846_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08171_ _00498_ _02100_ _02105_ _02109_ VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_37 _00953_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_15 _00722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 _01149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07122_ _01206_ VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_59 _01368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07053_ _01054_ Qset\[2\]\[13\] _01128_ VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07955_ _06279_ _01982_ _01960_ VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__a21o_1
X_06906_ _01023_ _01028_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__nand2_2
X_07886_ result_reg_Rshift\[15\] _01603_ _01601_ _01935_ VGND VGND VPWR VPWR _01936_
+ sky130_fd_sc_hd__o211a_1
X_09625_ _03532_ _03533_ VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__nand2_1
X_06837_ _00956_ _00961_ _00608_ VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__mux2_1
X_06768_ _00890_ _00709_ _00603_ _00895_ VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_87_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09556_ _03463_ _03464_ VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__nand2_1
X_06699_ _00574_ VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__inv_2
X_09487_ _03394_ _03396_ VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__nand2_1
X_08507_ _02311_ _02412_ _02139_ _02419_ _02426_ VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__o221ai_4
X_08438_ Qset\[0\]\[9\] VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08369_ _02248_ _02292_ _02254_ _02293_ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__o211ai_1
X_11380_ _05281_ _05254_ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__nand2_1
X_10400_ _04305_ _03768_ _00589_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__a21o_1
X_10331_ _04236_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10262_ _04166_ _04168_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__nand2_1
X_12001_ _04093_ _05749_ _04086_ _05745_ _05837_ VGND VGND VPWR VPWR _05838_ sky130_fd_sc_hd__a221o_1
X_10193_ _04052_ _04099_ VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__or2_1
X_12903_ clknet_leaf_16_clk _00346_ VGND VGND VPWR VPWR result_reg_and\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_88_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12834_ clknet_leaf_7_clk _00277_ VGND VGND VPWR VPWR result_reg_mul\[1\] sky130_fd_sc_hd__dfxtp_1
X_12765_ clknet_leaf_40_clk _00208_ VGND VGND VPWR VPWR H\[0\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_11716_ _05476_ VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12696_ clknet_leaf_36_clk _00146_ VGND VGND VPWR VPWR Oset\[0\]\[10\] sky130_fd_sc_hd__dfxtp_1
Xinput13 data_in[6] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
XFILLER_0_83_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11647_ _05545_ _05546_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput35 rst VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_2
Xinput24 instruction_in[16] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_2
X_11578_ _05477_ _05357_ _05478_ VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__nand3_1
XFILLER_0_52_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10529_ _04433_ _04434_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07740_ _01796_ result_reg_mac\[8\] _01570_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07671_ _01728_ _01663_ _01729_ _01730_ VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06622_ result_reg_Lshift\[2\] VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__inv_2
X_09410_ _03318_ _03319_ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09341_ _02908_ _02907_ _03251_ VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__a21oi_2
X_06553_ _00668_ Qset\[0\]\[0\] _00687_ VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__mux2_1
X_06484_ _00603_ VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__inv_2
X_09272_ _03150_ _03182_ VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08223_ _02151_ _02152_ _02147_ _02153_ VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__a211o_1
XFILLER_0_105_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08154_ _00547_ _02096_ current_state\[6\] VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07105_ _01189_ VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08085_ _01650_ H\[1\]\[1\] _02057_ VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__mux2_1
X_07036_ _01134_ VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08987_ _02619_ _02895_ VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__nand2_1
X_07938_ _01969_ VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07869_ _01919_ VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09608_ _03514_ _03509_ _03510_ VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__nand3_1
X_10880_ _04780_ _04783_ VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09539_ _03291_ _03448_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12550_ _01004_ Qset\[3\]\[11\] _06233_ VGND VGND VPWR VPWR _06246_ sky130_fd_sc_hd__mux2_1
X_12481_ _06181_ _06133_ _06149_ _06106_ VGND VGND VPWR VPWR _06206_ sky130_fd_sc_hd__a31oi_1
X_11501_ _05400_ _05401_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__nand2_1
X_11432_ _00585_ _02489_ _05332_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11363_ _05263_ _05262_ VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11294_ _05194_ _05193_ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10314_ _04218_ _04220_ VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__nand2_1
X_10245_ _04138_ _04140_ _04151_ VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__o21ai_1
X_10176_ _02523_ Oset\[2\]\[15\] VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_45_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12817_ clknet_leaf_10_clk _00260_ VGND VGND VPWR VPWR result_reg_sub\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12748_ clknet_leaf_37_clk _00191_ VGND VGND VPWR VPWR H\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12679_ clknet_leaf_1_clk _00129_ VGND VGND VPWR VPWR LC\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09890_ H\[3\]\[8\] _03793_ _03795_ _03796_ VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__a211o_1
X_08910_ _02619_ _02821_ VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__nand2_1
X_08841_ _02581_ Qset\[2\]\[2\] VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08772_ _02685_ _02192_ VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__nand2_1
X_07723_ _01613_ _01765_ _01780_ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__a21o_2
X_07654_ _01714_ result_reg_mac\[4\] _01570_ VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06605_ result_reg_or\[2\] VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__inv_2
X_07585_ result_reg_mac\[1\] _01541_ _01606_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06536_ R2\[1\] VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__inv_2
X_09324_ _02910_ _02912_ VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__nand2_1
X_06467_ _00575_ _00596_ _00601_ VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09255_ _03165_ VGND VGND VPWR VPWR _03166_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08206_ _02134_ _02135_ _02136_ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__nand3_1
XFILLER_0_28_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06398_ _00532_ VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09186_ _03093_ _03096_ VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08137_ H\[0\]\[10\] _01839_ _02074_ VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08068_ _01839_ H\[2\]\[10\] _02037_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__mux2_1
X_07019_ _01080_ Qset\[1\]\[14\] _01108_ VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__mux2_1
X_10030_ _03936_ _03878_ _03883_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_59_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11981_ _04891_ _05744_ _04107_ _05766_ _05820_ VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__a221o_2
X_10932_ _03764_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10863_ _04766_ _04578_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_104_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12602_ clknet_leaf_34_clk _00052_ VGND VGND VPWR VPWR Qset\[1\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_10794_ _04649_ _04697_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12533_ _06237_ VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12464_ _06098_ _06187_ _06192_ _06138_ _06193_ VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11415_ result_reg_add\[13\] _02648_ _05134_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__o21ai_1
X_12395_ _06126_ _00547_ VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__nand2_1
X_11346_ _05247_ VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13016_ clknet_leaf_43_clk _00459_ VGND VGND VPWR VPWR Qset\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11277_ _04929_ _05178_ VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__nor2_1
X_10228_ _04131_ _04133_ _04134_ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__o21bai_1
X_10159_ _04059_ _04065_ _01155_ _03095_ VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07370_ _00985_ _01266_ _01299_ _01443_ VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06321_ LC\[8\] VGND VGND VPWR VPWR _06282_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09040_ _02950_ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__inv_2
X_09942_ _03848_ _02723_ VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09873_ _03776_ _03777_ _03778_ _03779_ VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__o22a_2
X_08824_ _02686_ VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__inv_2
X_08755_ _02579_ Oset\[1\]\[1\] VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__nand2_1
X_07706_ _00901_ _01608_ _01600_ _01763_ VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_56_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ _02599_ _00005_ _02600_ VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__nand3_2
X_07637_ result_reg_not\[3\] _01633_ _01698_ VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__a21o_1
X_07568_ result_reg_Lshift\[1\] _01608_ _01600_ _01631_ VGND VGND VPWR VPWR _01632_
+ sky130_fd_sc_hd__a211o_1
X_06519_ _00632_ _00653_ VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__nor2_8
XFILLER_0_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09307_ _03217_ _03185_ VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_615 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07499_ _01170_ _01561_ VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09238_ _03114_ _03146_ VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09169_ _02619_ _03079_ VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11200_ _05089_ _05102_ VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__xor2_1
X_12180_ _03162_ _02998_ _05892_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__a21oi_1
X_11131_ _05032_ _05030_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11062_ _04881_ _02463_ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__nor2_1
X_10013_ _03918_ _03903_ VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11964_ _05766_ _02118_ _05792_ _05806_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__a31o_1
XFILLER_0_98_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11895_ _01158_ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__clkbuf_4
X_10915_ _04817_ _04818_ _04814_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__nand3_1
XFILLER_0_73_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10846_ _04727_ _04749_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10777_ _03759_ Oset\[0\]\[11\] VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__nor2_1
X_12516_ net70 _06220_ _06221_ _06227_ VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__o211a_1
X_12447_ _06123_ _06128_ _06256_ _06267_ _06134_ VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__a311o_1
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12378_ _06097_ CMD_logic_shift_right _04827_ _06121_ VGND VGND VPWR VPWR _00415_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11329_ _05114_ _05230_ VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__nand2_1
X_06870_ _00993_ _00615_ VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08540_ _02454_ _02457_ VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_53_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08471_ _02327_ _02391_ VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__nand2_1
X_07422_ result_reg_not\[14\] _01492_ _01168_ VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07353_ _01427_ _01255_ VGND VGND VPWR VPWR _01428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07284_ _01359_ _01245_ _01362_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__a21o_1
X_06304_ _06267_ _06261_ VGND VGND VPWR VPWR _06268_ sky130_fd_sc_hd__or2_1
X_09023_ _02926_ _02934_ _02540_ VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_92_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09925_ _03831_ _02573_ _00588_ VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__a21oi_1
X_09856_ _03760_ H\[3\]\[8\] _03761_ _03762_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_5_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ _02714_ _02720_ _01154_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__nand3_1
XFILLER_0_99_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _03693_ _03694_ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__or2_1
X_06999_ _00809_ Qset\[1\]\[4\] _01109_ VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__mux2_1
X_08738_ _02652_ VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__inv_2
XANTENNA_105 _01870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_116 _02474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_149 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_127 _05298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_138 _06218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08669_ _00005_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__buf_4
XFILLER_0_95_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10700_ _04603_ _04604_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11680_ _05578_ _05579_ VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_101_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10631_ _03899_ _04495_ VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__nor2_1
X_10562_ _04266_ _04466_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__nor2_1
X_12301_ _05766_ _03131_ _00669_ _02126_ _03144_ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__o221a_1
X_12232_ result_reg_or\[13\] _05960_ _06019_ _06021_ _02101_ VGND VGND VPWR VPWR _00369_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10493_ _04339_ _04398_ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__nand2_1
X_12163_ _02711_ _02661_ VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__nand2_1
X_12094_ _05907_ _03328_ _03128_ _05894_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__o31ai_1
X_11114_ _04766_ _04901_ _04904_ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__o21a_1
X_11045_ _04946_ _04920_ VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12996_ clknet_leaf_0_clk _00439_ VGND VGND VPWR VPWR R1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11947_ _05788_ _05790_ _05791_ VGND VGND VPWR VPWR _05792_ sky130_fd_sc_hd__and3_2
XFILLER_0_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11878_ _05732_ VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__inv_2
X_10829_ _04105_ _02413_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07971_ _01962_ _06283_ _01964_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__a21o_1
X_06922_ _01043_ _01034_ _00534_ VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__mux2_1
X_09710_ _03506_ _03304_ VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__nand2_1
X_06853_ _00974_ _00655_ _00657_ _00977_ _00666_ VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__a221o_1
X_09641_ _03548_ _03544_ VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06784_ result_reg_mul\[8\] VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09572_ _02611_ _02296_ _02584_ _03480_ VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_38_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08523_ _02438_ _02441_ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08454_ _02372_ _02373_ _02374_ _02375_ VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__a211o_1
XFILLER_0_92_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07405_ _01185_ _01032_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__nand2_1
X_08385_ _02309_ net60 _02170_ VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07336_ _00939_ _01208_ _01190_ _01411_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07267_ result_reg_mac\[5\] _01215_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__nor2_1
X_09006_ _02592_ Oset\[3\]\[3\] VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__nand2_1
X_07198_ result_reg_not\[2\] _01280_ _01168_ VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09908_ Qset\[3\]\[8\] _03136_ VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__nor2_1
X_09839_ _03745_ VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__buf_6
X_12850_ clknet_leaf_20_clk _00293_ VGND VGND VPWR VPWR result_reg_mac\[1\] sky130_fd_sc_hd__dfxtp_1
X_11801_ _05679_ VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__inv_2
X_12781_ clknet_leaf_24_clk _00224_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_1_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11732_ _05630_ VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11663_ _03790_ _03076_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__nand2_1
X_10614_ _04518_ _03951_ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__nand2_1
X_11594_ _05335_ _02510_ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10545_ _04320_ _03411_ VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__nand2_1
X_10476_ _04380_ _04378_ _04379_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_32_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12215_ _03874_ _01666_ _06007_ _01243_ _05928_ VGND VGND VPWR VPWR _06008_ sky130_fd_sc_hd__a221o_1
X_12146_ _05506_ _00524_ _05836_ _05873_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12077_ _01282_ _05873_ _05891_ _05893_ _02650_ VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__a221oi_1
X_11028_ _04747_ _04929_ _04930_ VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12979_ clknet_leaf_2_clk _00422_ VGND VGND VPWR VPWR CMD_set sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_27 _00859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_16 _00742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08170_ _02102_ _02103_ net42 VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_38 _00953_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07121_ _00559_ _01198_ VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__nand2_2
XANTENNA_49 _01150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07052_ _01142_ VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07954_ _06277_ LC\[5\] VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07885_ _01716_ _01103_ VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__nand2_1
X_06905_ _01024_ _00654_ _00656_ _01027_ _00665_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__a221o_1
X_06836_ _00957_ _00960_ _00732_ VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__mux2_1
X_09624_ _03374_ _03375_ _03376_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__a21boi_1
X_06767_ _00892_ _00743_ _00893_ _00894_ VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__a31o_1
X_09555_ _02963_ _02895_ VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06698_ _00557_ _00631_ _00634_ _00827_ VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__or4_1
X_09486_ _03395_ VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__inv_2
X_08506_ _02422_ _02425_ _01553_ VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__a21o_2
X_08437_ _02356_ Qset\[3\]\[9\] _02347_ _02358_ VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__a211o_1
XFILLER_0_92_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08368_ _02248_ Qset\[1\]\[6\] VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07319_ _01395_ result_reg_mul\[8\] _01263_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_83_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08299_ _02141_ Oset\[1\]\[3\] VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10330_ _04235_ _04236_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__nand2_1
X_10261_ _03959_ _04167_ _04164_ VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__o21ai_1
X_12000_ _00591_ _05836_ VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__nor2_1
X_10192_ _04075_ _04097_ _04098_ VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_92_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12902_ clknet_leaf_15_clk _00345_ VGND VGND VPWR VPWR result_reg_and\[5\] sky130_fd_sc_hd__dfxtp_2
X_12833_ clknet_leaf_2_clk _00276_ VGND VGND VPWR VPWR result_reg_mul\[0\] sky130_fd_sc_hd__dfxtp_2
X_12764_ clknet_leaf_37_clk _00207_ VGND VGND VPWR VPWR H\[0\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11715_ _05613_ _05614_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12695_ clknet_leaf_40_clk _00145_ VGND VGND VPWR VPWR Oset\[0\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11646_ _05453_ _05449_ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput14 data_in[7] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
Xinput25 instruction_in[17] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_2
X_11577_ _05471_ _02160_ _05472_ VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__nand3_1
XFILLER_0_52_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10528_ _04432_ _04406_ _04412_ VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_12_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10459_ _04363_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12129_ _05907_ _04847_ _04891_ _05878_ VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__o31ai_1
X_07670_ result_reg_mul\[5\] _01688_ _01667_ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_48_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06621_ _00643_ VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__buf_2
X_09340_ _02823_ _03241_ VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__nor2_1
X_06552_ _00686_ VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__buf_6
XFILLER_0_87_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09271_ _03178_ _03180_ _03181_ VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__a21oi_1
X_06483_ net1 _00600_ _00617_ VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08222_ H\[3\]\[0\] _02151_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__nor2_1
X_08153_ _00556_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__buf_4
XFILLER_0_43_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07104_ _01185_ _01188_ _01181_ VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__or3b_1
XFILLER_0_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08084_ _02058_ VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07035_ _00809_ Qset\[2\]\[4\] _01129_ VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08986_ _02685_ _02192_ _02897_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_89_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07937_ _01968_ LC\[1\] _01964_ VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__mux2_1
X_07868_ _01918_ H\[3\]\[14\] _01628_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__mux2_1
X_06819_ _00939_ _00709_ _00603_ _00944_ VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__o211a_1
X_07799_ _00989_ _01574_ _01850_ _01852_ _01569_ VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__a221o_1
X_09607_ _03511_ _03515_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09538_ _03446_ _03447_ VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__or2b_2
XFILLER_0_93_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09469_ _03378_ _03274_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__nand2_1
X_11500_ _05288_ _05280_ _05399_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__a21o_1
X_12480_ _06205_ VGND VGND VPWR VPWR _00433_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11431_ _03770_ _05324_ _01156_ _05331_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__o211a_1
X_11362_ _05262_ _05263_ VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10313_ _04213_ _04219_ _04214_ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11293_ _05193_ _05194_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__or2_1
X_10244_ _04142_ _04143_ _04150_ VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__nand3_2
X_10175_ _02529_ Oset\[3\]\[15\] _02535_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12816_ clknet_leaf_10_clk _00259_ VGND VGND VPWR VPWR result_reg_add\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_45_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12747_ clknet_leaf_41_clk _00190_ VGND VGND VPWR VPWR H\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12678_ clknet_leaf_0_clk _00128_ VGND VGND VPWR VPWR LC\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11629_ _05431_ _05429_ _05527_ _03048_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08840_ _00635_ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08771_ _02684_ _01551_ VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__nand2_1
X_07722_ _00880_ _01570_ _01779_ VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__a21oi_1
X_07653_ _01594_ _01707_ _01713_ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__o21ai_1
X_06604_ net9 _00696_ _00736_ VGND VGND VPWR VPWR _00737_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07584_ _01639_ _01569_ _01640_ _01570_ _01647_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__a311o_1
XFILLER_0_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09323_ _03229_ _03232_ _03233_ VGND VGND VPWR VPWR _03234_ sky130_fd_sc_hd__nand3_1
XFILLER_0_75_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06535_ R0\[1\] VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__inv_2
X_06466_ _00600_ VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09254_ _02562_ Oset\[1\]\[4\] VGND VGND VPWR VPWR _03165_ sky130_fd_sc_hd__nand2_1
X_09185_ _03095_ VGND VGND VPWR VPWR _03096_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08205_ Qset\[1\]\[0\] _02131_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06397_ _00528_ _00531_ VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__nor2_2
X_08136_ _02085_ VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08067_ _02048_ VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__clkbuf_1
X_07018_ _01123_ VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__clkbuf_1
X_08969_ _02875_ _02877_ _02880_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__o21ai_4
X_11980_ _02139_ _04886_ VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__nor2_1
X_10931_ H\[2\]\[12\] H\[3\]\[12\] _04283_ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10862_ _04074_ _03421_ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_104_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10793_ _04695_ _04696_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__xor2_2
XFILLER_0_38_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12601_ clknet_leaf_35_clk _00051_ VGND VGND VPWR VPWR Qset\[1\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12532_ _00759_ Qset\[3\]\[2\] _06234_ VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12463_ _06123_ _06112_ _06116_ _06266_ VGND VGND VPWR VPWR _06193_ sky130_fd_sc_hd__a31o_1
X_11414_ _05312_ _05314_ _05313_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_50_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12394_ _06104_ _06129_ _06122_ net25 _06135_ VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_104_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11345_ _05245_ _05246_ VGND VGND VPWR VPWR _05247_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11276_ _04690_ _04555_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_72_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13015_ clknet_leaf_44_clk _00458_ VGND VGND VPWR VPWR Qset\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_10227_ _03205_ _04110_ VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10158_ _04064_ _02552_ VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10089_ _03994_ _03995_ VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06320_ LC\[7\] _06280_ VGND VGND VPWR VPWR _06281_ sky130_fd_sc_hd__and2b_1
XFILLER_0_45_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09941_ _03841_ _01156_ _03847_ VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__nand3_1
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09872_ Qset\[1\]\[8\] _03773_ _03004_ VGND VGND VPWR VPWR _03779_ sky130_fd_sc_hd__o21ai_1
X_08823_ _02736_ _02621_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__or2_1
X_08754_ _02580_ Oset\[0\]\[1\] VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__nand2_1
X_07705_ result_reg_Rshift\[7\] _01608_ VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_56_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08685_ _02585_ Oset\[3\]\[0\] VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__nand2_1
X_07636_ result_reg_Rshift\[3\] _01672_ _01607_ _01697_ VGND VGND VPWR VPWR _01698_
+ sky130_fd_sc_hd__o211a_1
X_07567_ _00690_ _01608_ VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06518_ _00550_ VGND VGND VPWR VPWR _00653_ sky130_fd_sc_hd__inv_2
X_09306_ _03187_ _03183_ VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__nand2_1
X_07498_ _01557_ net1 _01558_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09237_ _03114_ _03147_ VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_35_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06449_ _00583_ VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09168_ _03051_ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__inv_2
X_08119_ H\[0\]\[1\] _01650_ _02075_ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__mux2_1
X_09099_ _03008_ _03009_ VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__nand2_1
X_11130_ _05030_ _05032_ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__or2_1
X_11061_ _02163_ _04963_ _02713_ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__o21ai_1
X_10012_ _03903_ _03918_ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11963_ _02118_ _05805_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11894_ _00590_ VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__clkbuf_4
X_10914_ _04792_ _02160_ _04793_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_27_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10845_ _04556_ _04745_ _04748_ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10776_ _03498_ Oset\[2\]\[11\] _03345_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12515_ _06219_ _00500_ VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__nand2_1
X_12446_ _06142_ _06178_ _06147_ _06106_ VGND VGND VPWR VPWR _06179_ sky130_fd_sc_hd__a31oi_1
X_12377_ _06120_ _06097_ VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__nand2_1
X_11328_ _05058_ _05110_ VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11259_ _04855_ Qset\[0\]\[13\] _04862_ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08470_ Qset\[0\]\[10\] VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__inv_2
X_07421_ result_reg_Lshift\[14\] result_reg_Rshift\[14\] _01165_ VGND VGND VPWR VPWR
+ _01492_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07352_ _00956_ _01426_ _01182_ VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06303_ _06266_ VGND VGND VPWR VPWR _06267_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_61_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07283_ _00860_ _01266_ _01206_ _01361_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09022_ _02933_ _00580_ VGND VGND VPWR VPWR _02934_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09924_ _03135_ _03828_ _03830_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__o21ai_4
X_09855_ _03760_ _02346_ VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08806_ _02719_ _02551_ VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_69_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09786_ _03385_ _03546_ _03550_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__o21a_1
X_06998_ _01113_ VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__clkbuf_1
X_08737_ _02646_ _02649_ _02650_ _02651_ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__a211o_1
XANTENNA_106 _01890_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_128 _05693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 _02545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_139 _06218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08668_ _02582_ Qset\[2\]\[0\] VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__nand2_1
X_07619_ _01678_ _01549_ _01680_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08599_ H\[1\]\[15\] _02327_ VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__nor2_1
X_10630_ _04532_ _04534_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_101_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10561_ _04275_ VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__inv_2
X_12300_ _01148_ VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__clkbuf_4
X_10492_ _04397_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__inv_2
X_12231_ _06020_ _00524_ _05154_ _01666_ _05943_ VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__a221o_1
XFILLER_0_51_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12162_ result_reg_or\[0\] _05959_ _05962_ _05964_ _05940_ VGND VGND VPWR VPWR _00356_
+ sky130_fd_sc_hd__o221a_1
X_12093_ _05892_ VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__clkbuf_4
X_11113_ _05012_ _05015_ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__xor2_1
X_11044_ _04920_ _04946_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12995_ clknet_leaf_15_clk _00438_ VGND VGND VPWR VPWR R0\[1\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_56_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11946_ _03063_ _01158_ VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11877_ _05132_ _05133_ _05703_ _05731_ VGND VGND VPWR VPWR _05732_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10828_ _04731_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__inv_2
X_10759_ _04661_ _04459_ _04662_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_15_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12429_ net21 _06131_ VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_78_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07970_ im_reg\[8\] _01962_ VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__nor2_1
X_06921_ _01035_ _01036_ _00539_ VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06852_ result_reg_Rshift\[10\] _00753_ _00976_ VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09640_ _03544_ _03548_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__or2_1
X_06783_ result_reg_or\[8\] _00553_ result_reg_and\[8\] _00562_ _00603_ VGND VGND
+ VPWR VPWR _00910_ sky130_fd_sc_hd__o221a_1
X_09571_ _02611_ Oset\[3\]\[6\] VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_66_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08522_ _02364_ Oset\[1\]\[12\] _02378_ _02440_ VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__a211o_1
XFILLER_0_26_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08453_ _02373_ H\[2\]\[9\] VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07404_ result_reg_not\[13\] _01475_ _01167_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08384_ _02126_ _02295_ _02140_ _02302_ _02308_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__o221ai_4
X_07335_ _01407_ _01207_ _01261_ _01410_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07266_ _01344_ _01199_ _01190_ _01345_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__a211o_1
XFILLER_0_73_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09005_ _02581_ Oset\[2\]\[3\] VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07197_ result_reg_Lshift\[2\] result_reg_Rshift\[2\] _01165_ VGND VGND VPWR VPWR
+ _01280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09907_ _03754_ _03756_ _03813_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__nand3_1
X_09838_ _03050_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__clkbuf_4
X_09769_ _03529_ _03531_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__nand2_1
X_11800_ _03234_ _03276_ _05670_ _05678_ VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_38_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12780_ clknet_leaf_24_clk _00223_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dfxtp_1
X_11731_ _05628_ _02645_ _05629_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__o21ai_1
X_11662_ _04308_ _03110_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11593_ _05424_ _05421_ VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__nand2_1
X_10613_ _03950_ _03948_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10544_ _04241_ _04240_ _04324_ VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__nand3_1
X_10475_ _04378_ _04379_ _04380_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__a21bo_1
X_12214_ _04546_ _04483_ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_102_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12145_ _01499_ _05873_ _02115_ _05949_ VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__a211oi_1
X_12076_ _05892_ _05750_ _02760_ _05878_ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__o31a_1
X_11027_ _04607_ _04495_ _04745_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
X_12978_ clknet_leaf_7_clk _00421_ VGND VGND VPWR VPWR CMD_store sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11929_ _00591_ _02118_ VGND VGND VPWR VPWR _05776_ sky130_fd_sc_hd__nand2_1
XANTENNA_17 _00750_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 _00871_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 _00972_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07120_ _01203_ result_reg_mul\[0\] _01204_ VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07051_ _01029_ Qset\[2\]\[12\] _01128_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07953_ _01981_ VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__clkbuf_1
X_07884_ _01933_ result_reg_mac\[15\] _01540_ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__mux2_1
X_06904_ result_reg_Rshift\[12\] _00753_ _01026_ VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06835_ _00958_ _00959_ _00730_ VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__mux2_1
X_09623_ _03530_ _03531_ VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__nand2_1
X_06766_ result_reg_and\[7\] _00561_ _00552_ VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09554_ _03020_ _03462_ VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__nand2_1
X_06697_ shift.left CMD_logic_shift_right _00820_ _00826_ VGND VGND VPWR VPWR _00827_
+ sky130_fd_sc_hd__or4_1
X_09485_ _03192_ _03197_ _03191_ VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__a21oi_2
X_08505_ _02423_ _02373_ _02378_ _02424_ VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08436_ _02328_ _02357_ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__nor2_1
X_08367_ Qset\[0\]\[6\] VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07318_ result_reg_add\[8\] result_reg_sub\[8\] _01264_ VGND VGND VPWR VPWR _01395_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08298_ Oset\[0\]\[3\] VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07249_ result_reg_mac\[4\] _01215_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10260_ _03942_ _03924_ VGND VGND VPWR VPWR _04167_ sky130_fd_sc_hd__and2_1
X_10191_ _04074_ _02687_ _04096_ _02620_ VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12901_ clknet_leaf_16_clk _00344_ VGND VGND VPWR VPWR result_reg_and\[4\] sky130_fd_sc_hd__dfxtp_1
X_12832_ clknet_leaf_10_clk _00275_ VGND VGND VPWR VPWR result_reg_sub\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12763_ clknet_leaf_41_clk _00206_ VGND VGND VPWR VPWR H\[0\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11714_ _05612_ _05593_ _05594_ VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_83_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12694_ clknet_leaf_42_clk _00144_ VGND VGND VPWR VPWR Oset\[0\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11645_ _05541_ _05544_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__xor2_1
Xinput15 data_in[8] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dlymetal6s2s_1
X_11576_ _05473_ _00832_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput26 instruction_in[1] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_40_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10527_ _04413_ _04432_ VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10458_ _04340_ _04363_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_75_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10389_ _04294_ _00582_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__nand2_1
X_12128_ _01851_ _05873_ _02115_ _05935_ VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__a211oi_1
X_12059_ _05871_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__clkbuf_4
X_06620_ _00643_ VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_48_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06551_ _00679_ _00685_ VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__nand2_4
XFILLER_0_59_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06482_ result_reg_set\[0\] _00608_ _00601_ _00616_ VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09270_ _03107_ _03179_ VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08221_ H\[2\]\[0\] VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08152_ _02094_ _00578_ _00546_ VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__and3_2
XFILLER_0_55_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_9_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
X_07103_ _01171_ _00568_ VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__nor2_1
X_08083_ _01615_ H\[1\]\[0\] _02057_ VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07034_ _01133_ VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08985_ _02821_ VGND VGND VPWR VPWR _02897_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_89_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07936_ _01967_ R3\[1\] _01960_ VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__mux2_1
X_07867_ _01914_ _01917_ _01612_ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__mux2_1
X_06818_ _00941_ _00743_ _00942_ _00943_ VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__a31o_1
X_07798_ _01571_ _00551_ _01851_ _01588_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__o2bb2a_1
X_09606_ _03514_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__inv_2
X_06749_ _00872_ _00877_ VGND VGND VPWR VPWR _00878_ sky130_fd_sc_hd__nand2_4
X_09537_ _03445_ _03299_ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09468_ _03373_ _03377_ VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__nand2_1
X_08419_ Oset\[2\]\[8\] Oset\[3\]\[8\] _02261_ VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__mux2_1
X_09399_ _03307_ _03308_ VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__nand2_1
X_11430_ _00582_ _05329_ _05330_ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11361_ _04458_ _04924_ VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10312_ _04217_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11292_ _04944_ _04941_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__nand2_1
X_10243_ _04149_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__inv_2
X_10174_ _04078_ _04080_ _00581_ _02871_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12815_ clknet_leaf_10_clk _00258_ VGND VGND VPWR VPWR result_reg_add\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_45_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_4__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_12746_ clknet_leaf_41_clk _00189_ VGND VGND VPWR VPWR H\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12677_ clknet_leaf_0_clk _00127_ VGND VGND VPWR VPWR LC\[1\] sky130_fd_sc_hd__dfxtp_1
X_11628_ _05431_ _05429_ _05527_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11559_ _05459_ _05042_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08770_ _02676_ _02683_ VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__nand2_1
X_07721_ _01771_ _01541_ _01778_ _01612_ VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__a31o_1
XFILLER_0_26_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07652_ _00795_ _01574_ _01711_ _01712_ _01569_ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__a221o_1
X_06603_ _00734_ _00735_ VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__nand2_1
X_07583_ _01574_ _01645_ _01593_ _01646_ VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__o211a_1
X_06534_ R3\[1\] VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__inv_2
X_09322_ _03051_ VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06465_ _00599_ VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__buf_2
X_09253_ _02565_ _02253_ VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__nor2_1
X_06396_ _00530_ VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__inv_2
X_09184_ _01154_ _03094_ _02555_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__o21ai_2
X_08204_ _00003_ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08135_ H\[0\]\[9\] _01819_ _02075_ VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_555 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08066_ _01819_ H\[2\]\[9\] _02038_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07017_ _01054_ Qset\[1\]\[13\] _01108_ VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08968_ _02878_ _02727_ _02879_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__nand3_1
X_07919_ _01955_ VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__clkbuf_1
X_08899_ _02809_ _02811_ VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__nand2_1
X_10930_ _02446_ _04832_ _03764_ VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10861_ _03507_ _04050_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12600_ clknet_leaf_34_clk _00050_ VGND VGND VPWR VPWR Qset\[1\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_104_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10792_ _04468_ _04496_ _04470_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_81_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12531_ _06236_ VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12462_ _06191_ _06186_ VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11413_ _05312_ _05313_ _05314_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_50_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12393_ _06254_ _06257_ _06134_ VGND VGND VPWR VPWR _06135_ sky130_fd_sc_hd__o21bai_1
X_11344_ _05077_ _05074_ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11275_ _04747_ _04929_ _04932_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_72_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10226_ _04132_ VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__inv_2
X_13014_ clknet_leaf_46_clk _00457_ VGND VGND VPWR VPWR Qset\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_10157_ _04061_ _04063_ VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__nor2_2
X_10088_ _03993_ _03988_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12729_ clknet_leaf_32_clk _00172_ VGND VGND VPWR VPWR H\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09940_ _03846_ _03781_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09871_ _03759_ Qset\[0\]\[8\] VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08822_ _02687_ _02734_ VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__nand2_1
X_08753_ _02665_ _00005_ _02666_ VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__nand3_2
X_07704_ _01762_ VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08684_ _02581_ Oset\[2\]\[0\] VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__nand2_1
X_07635_ _01608_ _00779_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07566_ _01630_ VGND VGND VPWR VPWR _00094_ sky130_fd_sc_hd__clkbuf_1
X_06517_ result_reg_not\[0\] VGND VGND VPWR VPWR _00652_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09305_ _03215_ VGND VGND VPWR VPWR _03216_ sky130_fd_sc_hd__inv_2
X_07497_ result_reg_mul\[0\] _01549_ _01559_ _01561_ VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09236_ _03146_ VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06448_ shift.O VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06379_ _00515_ _00511_ VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__or2_1
X_09167_ _03077_ VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__inv_2
X_09098_ _02257_ _00583_ _02572_ VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__a21oi_1
X_08118_ _02076_ VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__clkbuf_1
X_08049_ _02039_ VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__clkbuf_1
X_11060_ _04045_ _04960_ _04962_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_101_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10011_ _03904_ _03914_ _03917_ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11962_ _03840_ _05744_ _03846_ _05745_ _05804_ VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__a221o_2
XFILLER_0_98_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11893_ _05741_ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10913_ _04794_ _00832_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_27_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10844_ _04746_ _04025_ _04747_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12514_ net69 _06220_ _06221_ _06226_ VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__o211a_1
X_10775_ Oset\[3\]\[11\] _03341_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12445_ _06174_ VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__inv_2
X_12376_ net22 net25 _06254_ _06256_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11327_ _05228_ _04196_ VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11258_ _04855_ Qset\[2\]\[13\] VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11189_ _04458_ _04691_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__nor2_1
X_10209_ _04111_ _04113_ _04114_ _04115_ VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_82_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07420_ _01491_ VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07351_ _00957_ _01425_ _01177_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06302_ current_state\[2\] VGND VGND VPWR VPWR _06266_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07282_ _00865_ _01202_ _01204_ _01360_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_61_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09021_ _02929_ _02932_ VGND VGND VPWR VPWR _02933_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09923_ _02567_ H\[1\]\[8\] _02560_ _03829_ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__a211o_1
X_09854_ _03004_ VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__clkbuf_4
X_08805_ _02716_ _02718_ VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_69_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09785_ _03687_ _03692_ VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__xor2_1
X_06997_ _00783_ Qset\[1\]\[3\] _01109_ VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__mux2_1
X_08736_ result_reg_add\[0\] _02648_ VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__nor2_1
XANTENNA_107 _01909_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_129 _05711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_118 _02545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08667_ _02581_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__buf_6
X_07618_ result_reg_mul\[3\] _01679_ _01561_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08598_ H\[0\]\[15\] VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_101_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07549_ _00652_ _01607_ _01609_ _01610_ _01613_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__o221a_1
XFILLER_0_63_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10560_ _04463_ _04464_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09219_ _03123_ _03129_ _01155_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__nand3_1
X_10491_ _04392_ _04396_ VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__nand2_1
X_12230_ _05147_ _04963_ VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12161_ _05904_ _05746_ _01243_ _05963_ _05874_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12092_ result_reg_and\[4\] _05894_ _05901_ _05906_ _02125_ VGND VGND VPWR VPWR _00344_
+ sky130_fd_sc_hd__o221a_1
X_11112_ _05013_ _04954_ _05014_ VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__o21ai_1
X_11043_ _04944_ _04945_ VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_24_Left_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12994_ clknet_leaf_7_clk _00437_ VGND VGND VPWR VPWR R0\[0\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_4_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11945_ _05789_ _00590_ VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11876_ result_reg_mac\[12\] _05703_ _05682_ VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10827_ _04105_ Oset\[1\]\[11\] VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__nand2_1
X_10758_ _04265_ _04461_ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12428_ _06102_ _01962_ VGND VGND VPWR VPWR _06163_ sky130_fd_sc_hd__nor2_1
X_10689_ _04591_ _04387_ _04386_ VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__nand3_1
XFILLER_0_35_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12359_ _06098_ VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06920_ result_reg_and\[13\] VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__inv_2
X_06851_ _00754_ _00975_ VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__nand2_1
X_06782_ result_reg_mul\[8\] _00535_ _00907_ _00908_ _00563_ VGND VGND VPWR VPWR _00909_
+ sky130_fd_sc_hd__a221o_1
X_09570_ _02586_ Oset\[1\]\[6\] _02584_ VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_66_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08521_ _02364_ _02439_ VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08452_ _02347_ VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__clkbuf_4
X_07403_ result_reg_Lshift\[13\] result_reg_Rshift\[13\] _01164_ VGND VGND VPWR VPWR
+ _01475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08383_ _02305_ _02307_ _01552_ VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__a21o_2
X_07334_ _00931_ _01204_ _01244_ _01409_ VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__a211o_1
XFILLER_0_73_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07265_ result_reg_or\[5\] _01199_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09004_ _02914_ _02915_ VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__nand2_1
X_07196_ _01279_ VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09906_ _03811_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09837_ _03604_ _03734_ _03743_ VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__nand3_1
X_09768_ _03605_ _03675_ VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ Qset\[0\]\[0\] _02632_ _02633_ VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11730_ _05628_ _00610_ _02650_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__a21oi_1
X_09699_ _03606_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11661_ _05366_ _05363_ _05365_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11592_ _05491_ _05482_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10612_ _04516_ VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10543_ _04447_ VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10474_ _03350_ _04110_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__nor2_1
X_12213_ _05958_ _06005_ VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__nand2_1
X_12144_ _05945_ _05946_ _05878_ _05948_ VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__and4_1
X_12075_ _00525_ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__clkbuf_4
X_11026_ _04494_ _04744_ VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__nand2_1
X_12977_ clknet_leaf_7_clk _00420_ VGND VGND VPWR VPWR CMD_load sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11928_ _00635_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__buf_4
X_11859_ _00856_ _05707_ _05710_ _05719_ VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__a211o_1
XFILLER_0_86_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_18 _00759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 _00878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07050_ _01141_ VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07952_ _01980_ LC\[4\] _01964_ VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__mux2_1
X_07883_ _01593_ _01925_ _01932_ VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__o21ai_1
X_06903_ _00754_ _01025_ VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__nand2_1
X_06834_ result_reg_add\[10\] VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__inv_2
X_09622_ _03519_ _03520_ _03524_ VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__nand3_1
X_09553_ _03458_ VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__inv_2
X_06765_ _00882_ _00745_ VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__or2_1
X_08504_ _02397_ H\[0\]\[11\] VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06696_ CMD_not _00545_ CMD_and _00825_ VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__or4_1
XFILLER_0_65_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09484_ _03392_ _03393_ VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__nand2_1
X_08435_ Qset\[2\]\[9\] VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08366_ _02248_ _02289_ _02250_ _02290_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_18_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07317_ _01393_ _01255_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08297_ _02151_ Oset\[2\]\[3\] _02224_ VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07248_ _01327_ _01271_ _01254_ _01328_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07179_ _01204_ VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__clkbuf_4
X_10190_ _04096_ _02687_ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__nand2_1
X_12900_ clknet_leaf_15_clk _00343_ VGND VGND VPWR VPWR result_reg_and\[3\] sky130_fd_sc_hd__dfxtp_2
X_12831_ clknet_leaf_9_clk _00274_ VGND VGND VPWR VPWR result_reg_sub\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12762_ clknet_leaf_43_clk _00205_ VGND VGND VPWR VPWR H\[0\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11713_ _05595_ _05612_ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__nand2_1
X_12693_ clknet_leaf_40_clk _00143_ VGND VGND VPWR VPWR Oset\[0\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11644_ _05542_ _05543_ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput16 data_in[9] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
X_11575_ _05357_ _05474_ _05475_ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__nand3b_2
XTAP_TAPCELL_ROW_12_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput27 instruction_in[2] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_40_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10526_ _00710_ _04308_ _04431_ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__o21ai_1
X_10457_ _04360_ _04362_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_75_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10388_ _04291_ _04293_ VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__nand2_2
X_12127_ _05888_ _05932_ _05878_ _05933_ _05934_ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__o2111a_1
X_12058_ _01200_ _05876_ _02550_ VGND VGND VPWR VPWR _05877_ sky130_fd_sc_hd__or3_1
X_11009_ _04910_ _04911_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_48_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06550_ _00684_ VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06481_ _00614_ _00615_ VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08220_ _02128_ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__buf_2
XFILLER_0_43_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08151_ CMD_store CMD_load _00597_ _02093_ VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07102_ _01186_ VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__buf_2
XFILLER_0_15_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08082_ _02056_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__buf_4
X_07033_ _00783_ Qset\[2\]\[3\] _01129_ VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08984_ _02822_ _02620_ _02895_ VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__nand3_1
X_07935_ _06273_ _01966_ VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__nand2_1
X_07866_ result_reg_not\[14\] _01600_ _01916_ VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09605_ _03512_ _03351_ _03513_ VGND VGND VPWR VPWR _03514_ sky130_fd_sc_hd__a21oi_2
X_06817_ result_reg_and\[9\] _00561_ _00552_ VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__o21ai_1
X_07797_ result_reg_and\[11\] VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__inv_2
X_06748_ _00873_ _00655_ _00657_ _00876_ _00666_ VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09536_ _03299_ _03445_ VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__nor2_1
X_09467_ _03374_ _03375_ _03376_ VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__nand3_1
X_08418_ _02337_ _02338_ _02339_ _02340_ VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__o22a_2
XFILLER_0_19_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06679_ _00809_ Qset\[0\]\[4\] _00687_ VGND VGND VPWR VPWR _00810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09398_ _02785_ _02895_ VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__nand2_1
X_08349_ _02241_ _02274_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11360_ _05094_ _05259_ _05261_ VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10311_ _04215_ _04217_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11291_ _05192_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__inv_2
X_10242_ _04146_ _04148_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__nand2_1
X_10173_ _02565_ _02500_ _04079_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_28_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12814_ clknet_leaf_9_clk _00257_ VGND VGND VPWR VPWR result_reg_add\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12745_ clknet_leaf_32_clk _00188_ VGND VGND VPWR VPWR H\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12676_ clknet_leaf_0_clk _00126_ VGND VGND VPWR VPWR LC\[0\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_7_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11627_ _05493_ _05526_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11558_ _05041_ _05028_ VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10509_ _04414_ VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__clkbuf_4
X_11489_ _05388_ _05389_ VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_12_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07720_ _00890_ _01574_ _01775_ _01777_ _01569_ VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07651_ _01571_ _00551_ _01323_ _01667_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__o2bb2a_1
X_07582_ _01574_ _00708_ VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__nand2_1
X_06602_ _00699_ VGND VGND VPWR VPWR _00735_ sky130_fd_sc_hd__clkbuf_4
X_06533_ _00630_ _00645_ _00651_ _00667_ VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__a31o_2
X_09321_ _03230_ _03231_ VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__nand2_1
X_06464_ _00595_ _00598_ VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09252_ _02162_ _03162_ _02542_ VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__o21ai_1
X_06395_ current_state\[5\] _00529_ VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__nor2_2
X_09183_ im_reg\[6\] VGND VGND VPWR VPWR _03094_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08203_ _02129_ Qset\[0\]\[0\] VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08134_ _02084_ VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08065_ _02047_ VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07016_ _01122_ VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__clkbuf_1
X_08967_ _02874_ Oset\[3\]\[3\] VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07918_ Oset\[2\]\[12\] _01473_ _01941_ VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__mux2_1
X_08898_ _02810_ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__inv_2
X_07849_ _01067_ _01057_ _01544_ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__mux2_1
X_10860_ _04580_ _04577_ _04579_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09519_ _03021_ Oset\[2\]\[5\] VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_104_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10791_ _04693_ _04694_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__nand2_2
XFILLER_0_93_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12530_ _00722_ Qset\[3\]\[1\] _06234_ VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12461_ _06189_ _06190_ VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11412_ _05128_ _05130_ _04876_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_50_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12392_ _06130_ _06133_ VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11343_ _05232_ _05244_ VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_89_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11274_ _04926_ _05158_ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_72_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10225_ _04130_ _04122_ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__nand2_1
X_13013_ clknet_leaf_48_clk _00456_ VGND VGND VPWR VPWR Qset\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_10156_ Oset\[1\]\[14\] _02523_ _02535_ _04062_ VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__o211a_1
X_10087_ _03988_ _03993_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10989_ _02163_ _04891_ _02542_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12728_ clknet_leaf_44_clk _00171_ VGND VGND VPWR VPWR H\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_12659_ clknet_leaf_26_clk _00109_ VGND VGND VPWR VPWR H\[3\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09870_ _03759_ Qset\[2\]\[8\] _03345_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__o21ai_1
X_08821_ _02734_ VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08752_ _02579_ Oset\[3\]\[1\] VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__nand2_1
X_07703_ _01761_ H\[3\]\[6\] _01629_ VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__mux2_1
X_08683_ _02596_ _02597_ _02539_ VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__nand3_1
X_07634_ _01695_ result_reg_mac\[3\] _01570_ VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07565_ _01615_ H\[3\]\[0\] _01629_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__mux2_1
X_07496_ _01560_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__buf_2
X_06516_ result_reg_mac\[0\] _00650_ VGND VGND VPWR VPWR _00651_ sky130_fd_sc_hd__or2b_1
XFILLER_0_75_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09304_ _03213_ _03189_ VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09235_ _03116_ _03145_ VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__nand2_1
X_06447_ _00581_ VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__buf_4
XFILLER_0_90_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06378_ next_PC\[8\] VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__inv_2
X_09166_ _03052_ _03076_ VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09097_ _03000_ _01154_ _03007_ VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__nand3_1
X_08117_ H\[0\]\[0\] _01615_ _02075_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__mux2_1
X_08048_ _01615_ H\[2\]\[0\] _02038_ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10010_ _03915_ _03916_ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__nand2_1
X_09999_ _03835_ _02785_ _03050_ VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__nand3_1
X_11961_ _01554_ _05803_ VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__nor2_1
X_10912_ _04795_ _04796_ _04815_ VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__nand3_2
X_11892_ _05742_ VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_55_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10843_ _04308_ _04555_ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10774_ _04677_ _00582_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12513_ next_PC\[4\] _06218_ VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12444_ _06169_ _06177_ _02116_ VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_97_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12375_ _06118_ _06102_ _02115_ _06119_ VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_62_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11326_ _03751_ _05207_ _05227_ VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11257_ Qset\[3\]\[13\] _04857_ _04859_ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__a21oi_1
X_11188_ _04658_ _04654_ _04653_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__a21oi_1
X_10208_ _04074_ _02687_ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__nand2_1
X_10139_ _02567_ H\[3\]\[13\] _04045_ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07350_ _00958_ _00959_ _01174_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__mux2_1
X_06301_ _06265_ VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07281_ result_reg_add\[6\] _01202_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09020_ _02930_ _02591_ _02931_ VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__nand3_1
XFILLER_0_103_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09922_ _02565_ _02350_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__nor2_1
X_09853_ _03759_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__buf_6
X_08804_ _02527_ _02179_ _00007_ _02717_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__o211ai_1
X_09784_ _03689_ _03691_ VGND VGND VPWR VPWR _03692_ sky130_fd_sc_hd__nand2_1
X_08735_ _00635_ VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_69_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06996_ _01112_ VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_108 _01914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08666_ _02580_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__buf_6
XANTENNA_119 _02840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07617_ _01548_ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__clkbuf_4
X_08597_ _02509_ _02512_ VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_52_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07548_ _01612_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_101_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07479_ _00538_ _01543_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__nand2_4
XFILLER_0_63_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09218_ _02161_ _03128_ _02713_ VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__o21ai_1
X_10490_ _04393_ _04394_ _04395_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__nand3_1
X_09149_ _02874_ Oset\[3\]\[7\] _02534_ _03059_ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__a211o_1
X_12160_ _02550_ _05876_ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11111_ _03652_ _04074_ _04901_ VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_102_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12091_ _05902_ _01243_ _05903_ _05904_ _05905_ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11042_ _04921_ _04922_ _04943_ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__nand3_1
XFILLER_0_98_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12993_ clknet_leaf_7_clk _00436_ VGND VGND VPWR VPWR Qim sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11944_ _03054_ _03056_ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11875_ _05730_ VGND VGND VPWR VPWR _00303_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10826_ _04729_ _02416_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10757_ _04461_ _04265_ VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10688_ _04574_ _04592_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__nand2_1
X_12427_ _06161_ _06162_ _02116_ VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12358_ _06104_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__inv_2
X_12289_ _06054_ VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__inv_2
X_11309_ _04995_ _05210_ VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06850_ result_reg_Lshift\[10\] VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06781_ result_reg_sub\[8\] _00540_ VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08520_ Oset\[0\]\[12\] VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_38_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08451_ _02364_ VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07402_ _01474_ VGND VGND VPWR VPWR _00086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08382_ _02260_ H\[3\]\[6\] _02306_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07333_ _01204_ _01408_ VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07264_ result_reg_and\[5\] _01299_ _01343_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09003_ _02912_ _02902_ _02909_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__nand3_1
XFILLER_0_60_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07195_ Oset\[3\]\[1\] _01278_ _01250_ VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09905_ _03757_ _03811_ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__nand2_1
X_09836_ _03729_ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__inv_2
X_06979_ _00650_ _01098_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__nor2_1
X_09767_ _03672_ _03674_ VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ Qset\[1\]\[0\] _02624_ _00001_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__a21o_1
X_09698_ _03514_ _03511_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08649_ _02563_ VGND VGND VPWR VPWR _02564_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11660_ _04690_ _05078_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__nand2_1
X_11591_ _05484_ _05490_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__nand2_1
X_10611_ _04514_ _04515_ VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10542_ _04336_ _04334_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12212_ _04552_ _04477_ _05907_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10473_ _04377_ _04373_ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__nand2_1
X_12143_ _05947_ _05338_ VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_9_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12074_ _05888_ _02817_ _02781_ _05890_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__o31a_1
X_11025_ _04690_ _03859_ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__nand2_1
X_12976_ clknet_leaf_7_clk _00419_ VGND VGND VPWR VPWR CMD_not sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_63_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ _05741_ VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11858_ _05706_ _03601_ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__nor2_1
X_11789_ result_reg_mul\[0\] _05670_ _02105_ _05671_ VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__o211a_1
XANTENNA_19 _00759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10809_ _03956_ _04712_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__or2b_1
XFILLER_0_15_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07951_ _00498_ _01962_ _01978_ _01979_ VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06902_ result_reg_Lshift\[12\] VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__inv_2
X_07882_ _01929_ _01572_ _01930_ _01568_ _01931_ VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__a311o_1
X_06833_ result_reg_sub\[10\] VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__inv_2
X_09621_ _03521_ _03523_ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__nand2_1
X_06764_ result_reg_sub\[7\] _00740_ _00891_ VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__o21ai_1
X_09552_ _03348_ _02286_ _03303_ VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__a21oi_1
X_08503_ H\[1\]\[11\] VGND VGND VPWR VPWR _02423_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06695_ _00592_ CMD_set VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09483_ _03391_ _03384_ VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__nand2_1
X_08434_ _02319_ VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_43_Left_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08365_ _02261_ Qset\[3\]\[6\] VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__nand2_1
X_07316_ _01390_ _01392_ _01182_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08296_ _02223_ _02143_ VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__nand2_1
X_07247_ result_reg_or\[4\] _01199_ VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07178_ result_reg_and\[1\] _01207_ _01261_ VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_52_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09819_ _00624_ _03652_ _03726_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__o21ai_2
X_12830_ clknet_leaf_8_clk _00273_ VGND VGND VPWR VPWR result_reg_sub\[13\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_61_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12761_ clknet_leaf_32_clk _00204_ VGND VGND VPWR VPWR H\[0\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_11712_ _00832_ _05611_ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__xor2_1
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12692_ clknet_leaf_44_clk _00142_ VGND VGND VPWR VPWR Oset\[0\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_11643_ _05447_ _05443_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11574_ _05471_ _00832_ _05472_ VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__nand3_1
Xinput17 instruction_in[0] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_12_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput28 instruction_in[3] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_40_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10525_ _01537_ _04417_ _04419_ _00556_ _04430_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__a311o_2
XPHY_EDGE_ROW_70_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10456_ _04361_ _04341_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_75_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12126_ _05881_ _04683_ _04735_ VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__or3_1
X_10387_ _03760_ Qset\[1\]\[9\] _03764_ _04292_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__a211o_1
X_12057_ _02601_ _02604_ VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11008_ _04025_ _04899_ _04909_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_48_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ clknet_leaf_2_clk _00402_ VGND VGND VPWR VPWR result_reg_set\[14\] sky130_fd_sc_hd__dfxtp_1
X_06480_ _00607_ VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__buf_2
XFILLER_0_47_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08150_ _02092_ CMD_addition VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07101_ _01185_ VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__inv_2
X_08081_ _02055_ _01627_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__nand2b_4
X_07032_ _01132_ VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08983_ _02893_ _02894_ VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__nand2_4
X_07934_ LC\[1\] LC\[0\] VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07865_ result_reg_Rshift\[14\] _01603_ _01601_ _01915_ VGND VGND VPWR VPWR _01916_
+ sky130_fd_sc_hd__o211a_1
X_09604_ _03316_ _03314_ VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__nor2_1
X_06816_ _00931_ _00744_ VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__or2_1
X_07796_ _01847_ _01663_ _01848_ _01849_ VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06747_ result_reg_Rshift\[6\] _00753_ _00875_ VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09535_ _03440_ _03444_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__nand2_1
X_06678_ _00664_ _00803_ _00808_ VGND VGND VPWR VPWR _00809_ sky130_fd_sc_hd__o21ai_4
X_09466_ _03362_ _03365_ _03369_ VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__nand3_1
XFILLER_0_65_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08417_ Qset\[1\]\[8\] _02260_ _02254_ VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09397_ _02963_ _02821_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__nand2_1
X_08348_ Oset\[2\]\[5\] VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__inv_2
X_08279_ H\[3\]\[2\] _02151_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__nor2_1
X_10310_ _03790_ _04216_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__nand2_1
X_11290_ _05190_ _05191_ VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__nand2_1
X_10241_ _04112_ _04147_ VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__nor2_1
X_10172_ _03157_ Qset\[3\]\[15\] _02535_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__a21oi_1
X_12813_ clknet_leaf_9_clk _00256_ VGND VGND VPWR VPWR result_reg_add\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_45_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12744_ clknet_leaf_45_clk _00187_ VGND VGND VPWR VPWR H\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12675_ clknet_leaf_30_clk _00125_ VGND VGND VPWR VPWR Oset\[2\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11626_ _05518_ _05525_ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11557_ _05456_ _05457_ VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10508_ _03023_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11488_ _05387_ _05381_ VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__nand2_1
X_10439_ _03859_ VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12109_ _05888_ _03767_ _03831_ _05919_ VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_88_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07650_ _01708_ _01585_ _01709_ _01710_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__a31o_1
X_06601_ _00726_ _00733_ _00608_ VGND VGND VPWR VPWR _00734_ sky130_fd_sc_hd__mux2_1
X_07581_ _00715_ _01577_ _01644_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__o21ai_1
X_06532_ _00652_ _00655_ _00657_ _00660_ _00666_ VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_48_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09320_ _03228_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09251_ _03159_ _03161_ VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__nand2_1
X_06463_ _00597_ CMD_load _00578_ VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08202_ _02130_ _00003_ _02132_ VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__nand3_1
XFILLER_0_90_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06394_ _00471_ VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__inv_2
X_09182_ _03086_ _01155_ _03092_ VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__nand3_1
XFILLER_0_16_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08133_ H\[0\]\[8\] _01801_ _02075_ VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__mux2_1
X_08064_ _01801_ H\[2\]\[8\] _02038_ VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07015_ _01029_ Qset\[1\]\[12\] _01108_ VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08966_ _02522_ Oset\[2\]\[3\] VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__nand2_1
X_08897_ _00681_ _01154_ _02555_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__o21ai_1
X_07917_ _01954_ VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__clkbuf_1
X_07848_ _01899_ VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__clkbuf_1
X_07779_ _01594_ _01826_ _01833_ VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__o21ai_1
X_09518_ Oset\[3\]\[5\] _03024_ _02837_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__a21oi_1
X_10790_ _04692_ _04665_ _04666_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_38_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09449_ _03354_ _03358_ VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__nand2_1
X_12460_ net23 _06257_ VGND VGND VPWR VPWR _06190_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11411_ _05310_ _05308_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__nand2_1
X_12391_ _06132_ _06105_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_50_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11342_ _05242_ _05243_ VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__and2b_1
XFILLER_0_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11273_ _00820_ _05158_ _05174_ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10224_ _04122_ _04130_ VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__nor2_1
X_13012_ clknet_leaf_48_clk _00455_ VGND VGND VPWR VPWR Qset\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_10155_ _02523_ _02486_ VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10086_ _03990_ _03992_ VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_58_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10988_ _04045_ _04888_ _04890_ VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__o21ai_4
X_12727_ clknet_leaf_49_clk _00170_ VGND VGND VPWR VPWR H\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_12658_ clknet_leaf_27_clk _00108_ VGND VGND VPWR VPWR H\[3\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_11609_ _00585_ _02513_ _05508_ VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
X_12589_ clknet_leaf_26_clk _00039_ VGND VGND VPWR VPWR Qset\[0\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08820_ _02732_ _02733_ VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__nand2_2
X_08751_ _02580_ Oset\[2\]\[1\] VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07702_ _01757_ _01760_ _01613_ VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__mux2_4
X_08682_ _02138_ _02161_ VGND VGND VPWR VPWR _02597_ sky130_fd_sc_hd__nand2_1
X_07633_ _01594_ _01685_ _01694_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07564_ _01628_ VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__clkbuf_8
X_06515_ _00649_ VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__dlymetal6s2s_1
X_07495_ _01557_ _01180_ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__nand2_2
XFILLER_0_63_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09303_ _03189_ _03213_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09234_ _03143_ _03144_ VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__nand2_4
X_06446_ _00580_ VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09165_ _03074_ _03075_ VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__nand2_4
XFILLER_0_8_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06377_ _00513_ _00475_ _00514_ next_PC\[7\] _00478_ VGND VGND VPWR VPWR _00021_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08116_ _02074_ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__clkbuf_8
X_09096_ _03003_ _03006_ _02551_ VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__nand3_1
XFILLER_0_31_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08047_ _02037_ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09998_ _03886_ _03891_ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__xnor2_1
X_08949_ _00729_ _02654_ _02753_ _02861_ VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__a211o_1
X_11960_ _03854_ VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10911_ _04814_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__inv_2
X_11891_ _00659_ _02115_ _05741_ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_55_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10842_ _04744_ VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10773_ _04674_ _04676_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12512_ net68 _06220_ _06221_ _06225_ VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__o211a_1
X_12443_ _06173_ _06176_ _06267_ VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12374_ _06102_ _04830_ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11325_ _05225_ _03751_ _05226_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__nand3_1
X_11256_ _05157_ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__buf_6
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11187_ _04281_ _04924_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__nor2_1
X_10207_ _04049_ _02620_ VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__nand2_1
X_10138_ _03135_ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__buf_4
X_10069_ _03974_ _03975_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07280_ result_reg_and\[6\] VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__inv_2
X_06300_ _06263_ _06264_ _06261_ VGND VGND VPWR VPWR _06265_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09921_ H\[2\]\[8\] H\[3\]\[8\] _02529_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__mux2_1
X_09852_ _03498_ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__buf_6
X_08803_ _02527_ Oset\[3\]\[1\] VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__nand2_1
X_09783_ _03545_ _03690_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__nand2_1
X_08734_ _02648_ VGND VGND VPWR VPWR _02649_ sky130_fd_sc_hd__buf_4
X_06995_ _00759_ Qset\[1\]\[2\] _01109_ VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 _01929_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08665_ _02579_ VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__inv_4
X_07616_ _00770_ _00762_ _01545_ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__mux2_1
X_08596_ _02491_ Oset\[1\]\[15\] _02444_ _02511_ VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_52_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07547_ _01611_ VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__buf_4
XFILLER_0_76_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07478_ _01542_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06429_ result_reg_mul\[0\] _00535_ _00543_ _00544_ _00563_ VGND VGND VPWR VPWR _00564_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09217_ _03125_ _03127_ VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_32_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09148_ _02561_ _02320_ VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09079_ _02582_ Qset\[2\]\[4\] VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__nand2_1
X_11110_ _04074_ _03506_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__nand2_1
X_12090_ _03015_ _03155_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__nor2_1
X_11041_ _04921_ _04922_ _04943_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12992_ clknet_leaf_2_clk _00435_ VGND VGND VPWR VPWR Qreg3 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11943_ _03072_ _05749_ VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11874_ _05707_ _04826_ _05729_ VGND VGND VPWR VPWR _05730_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10825_ _04105_ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__buf_4
XFILLER_0_94_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10756_ _04657_ _04659_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10687_ _04591_ VGND VGND VPWR VPWR _04592_ sky130_fd_sc_hd__inv_2
X_12426_ _06126_ CMD_loopjump VGND VGND VPWR VPWR _06162_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12357_ net22 net23 VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12288_ R3\[1\] _06055_ _06044_ _06057_ VGND VGND VPWR VPWR _00389_ sky130_fd_sc_hd__o211a_1
X_11308_ _04690_ _04982_ VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__nand2_1
X_11239_ _04303_ _05137_ _05138_ _05139_ _05140_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__o32a_2
XFILLER_0_93_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06780_ _00541_ _00906_ _00535_ VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_66_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08450_ H\[3\]\[9\] VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07401_ Oset\[3\]\[12\] _01473_ _01249_ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__mux2_1
X_08381_ _02261_ H\[2\]\[6\] _02250_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__o21a_1
X_07332_ result_reg_add\[9\] result_reg_sub\[9\] _01201_ VGND VGND VPWR VPWR _01408_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07263_ result_reg_mul\[5\] _01263_ _01245_ _01342_ VGND VGND VPWR VPWR _01343_ sky130_fd_sc_hd__a211o_1
X_07194_ _01161_ _01253_ _01274_ _01277_ VGND VGND VPWR VPWR _01278_ sky130_fd_sc_hd__a22o_4
XFILLER_0_60_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09002_ _02910_ _02913_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09904_ _00624_ _03790_ _03810_ VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_6_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09835_ _03742_ VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__inv_2
X_06978_ net7 _00699_ _00839_ _01097_ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__o211a_1
X_09766_ _03667_ _03668_ _03673_ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__nand3_1
XFILLER_0_68_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08717_ _02624_ VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__inv_2
X_09697_ _03528_ _03530_ _03531_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08648_ H\[1\]\[0\] _02562_ VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__nand2_1
X_08579_ _02494_ _02491_ _02444_ _02495_ VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__a211o_1
X_11590_ _05483_ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10610_ _04512_ _04449_ _04453_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__nand3_1
XFILLER_0_36_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10541_ _04446_ VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12211_ result_reg_or\[9\] _05960_ _06002_ _06004_ _02101_ VGND VGND VPWR VPWR _00365_
+ sky130_fd_sc_hd__o221a_1
X_10472_ _04373_ _04377_ VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12142_ _01578_ _04071_ VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_9_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12073_ _01200_ _05889_ _02807_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__or3_1
X_11024_ _04748_ _04727_ _04556_ _04745_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__o2bb2a_1
X_12975_ clknet_leaf_7_clk _00418_ VGND VGND VPWR VPWR CMD_or sky130_fd_sc_hd__dfxtp_1
X_11926_ _05773_ VGND VGND VPWR VPWR _00311_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11857_ _05718_ VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__inv_2
X_11788_ _02621_ _05670_ VGND VGND VPWR VPWR _05671_ sky130_fd_sc_hd__nand2_1
X_10808_ _03955_ _03951_ VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10739_ _00959_ _02654_ _02753_ _04643_ VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__a211o_1
XFILLER_0_82_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12409_ _06147_ _06257_ _06100_ _06122_ _06253_ VGND VGND VPWR VPWR _06148_ sky130_fd_sc_hd__a41o_1
XFILLER_0_2_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07950_ _06277_ _01962_ VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06901_ result_reg_not\[12\] VGND VGND VPWR VPWR _01024_ sky130_fd_sc_hd__inv_2
X_07881_ result_reg_or\[15\] _01595_ VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__nor2_1
X_06832_ result_reg_mul\[10\] VGND VGND VPWR VPWR _00957_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09620_ _03527_ _03528_ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__nand2_1
X_06763_ _00540_ _00884_ _00534_ VGND VGND VPWR VPWR _00891_ sky130_fd_sc_hd__a21oi_1
X_09551_ _03459_ _03301_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__nand2_1
X_08502_ _02420_ _02373_ _02374_ _02421_ VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__a211o_1
X_06694_ _00557_ _00631_ _00823_ VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__or3_1
X_09482_ _03384_ _03391_ VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08433_ _02355_ VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08364_ Qset\[2\]\[6\] VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07315_ _00911_ _01391_ _01177_ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08295_ _02131_ Oset\[3\]\[3\] VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07246_ _01323_ _01245_ _01326_ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07177_ _00551_ _01243_ VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__nand2_4
X_09818_ _01537_ _03711_ _03713_ _00549_ _03725_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__a311o_2
X_09749_ _03619_ _03624_ _03610_ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__nand3_1
X_12760_ clknet_leaf_45_clk _00203_ VGND VGND VPWR VPWR H\[0\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11711_ _04830_ _05517_ _05610_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__o21ai_1
X_12691_ clknet_leaf_45_clk _00141_ VGND VGND VPWR VPWR Oset\[0\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11642_ _05517_ _04925_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__nand2_1
Xinput18 instruction_in[10] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
X_11573_ _05473_ _02160_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10524_ _04424_ _04429_ _01537_ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__a21oi_1
Xinput29 instruction_in[4] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_1
X_10455_ _04358_ _04359_ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12125_ _00525_ _04741_ _04677_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__or3_1
X_10386_ _03760_ _02360_ VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__nor2_1
X_12056_ _05874_ _05746_ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11007_ _04025_ _04899_ _04909_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12958_ clknet_leaf_1_clk _00401_ VGND VGND VPWR VPWR result_reg_set\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12889_ clknet_leaf_24_clk _00332_ VGND VGND VPWR VPWR result_reg_Rshift\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11909_ _01158_ _02719_ _02730_ _05749_ VGND VGND VPWR VPWR _05758_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07100_ _01179_ CMD_load _01184_ VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__and3_2
X_08080_ _01619_ _01622_ VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__nand2_1
X_07031_ _00759_ Qset\[2\]\[2\] _01129_ VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08982_ _00586_ R2\[1\] VGND VGND VPWR VPWR _02894_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07933_ _01961_ _01964_ _01965_ VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__o21ai_1
X_07864_ _01716_ _01076_ VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__nand2_1
X_06815_ result_reg_sub\[9\] _00740_ _00940_ VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__o21ai_1
X_09603_ _03314_ _03316_ VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__nand2_1
X_07795_ result_reg_mul\[11\] _01688_ _01589_ VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06746_ _00754_ _00874_ VGND VGND VPWR VPWR _00875_ sky130_fd_sc_hd__nand2_1
X_09534_ _03441_ _03442_ _03443_ VGND VGND VPWR VPWR _03444_ sky130_fd_sc_hd__nand3_1
X_06677_ _00804_ _00655_ _00657_ _00807_ _00666_ VGND VGND VPWR VPWR _00808_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09465_ _03275_ VGND VGND VPWR VPWR _03375_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08416_ _02319_ Qset\[0\]\[8\] VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09396_ _03305_ VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08347_ _02269_ _02272_ VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08278_ H\[2\]\[2\] VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__inv_2
X_07229_ net10 _01187_ _01254_ _01310_ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10240_ _04109_ _02620_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__nand2_2
X_10171_ _03136_ _04076_ _04077_ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_44_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12812_ clknet_leaf_10_clk _00255_ VGND VGND VPWR VPWR result_reg_add\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_45_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12743_ clknet_leaf_49_clk _00186_ VGND VGND VPWR VPWR H\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12674_ clknet_leaf_26_clk _00124_ VGND VGND VPWR VPWR Oset\[2\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_11625_ _05519_ _05524_ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__xor2_1
X_11556_ _05196_ _05190_ _05455_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10507_ _04406_ _04412_ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11487_ _05381_ _05387_ VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10438_ _04018_ _04014_ VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__and2_1
X_10369_ _04273_ _04274_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__nand2_1
X_12108_ _05892_ _03780_ _03819_ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__or3_1
X_12039_ result_reg_Rshift\[11\] _05847_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_88_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06600_ _00727_ _00731_ _00732_ VGND VGND VPWR VPWR _00733_ sky130_fd_sc_hd__mux2_1
X_07580_ _01641_ _01585_ _01642_ _01643_ VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__a31o_1
X_06531_ _00665_ VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09250_ _03136_ Qset\[2\]\[4\] _03160_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06462_ CMD_set _00545_ VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08201_ Qset\[3\]\[0\] _02131_ VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__nand2_1
X_06393_ CMD_multiplication VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__inv_2
X_09181_ _03091_ _02552_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08132_ _02083_ VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__clkbuf_1
X_08063_ _02046_ VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07014_ _01121_ VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08965_ _02876_ _02534_ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__nand2_1
X_07916_ Oset\[2\]\[11\] _01455_ _01941_ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__mux2_1
X_08896_ _02797_ _02808_ _01155_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__nand3_1
X_07847_ _01898_ H\[3\]\[13\] _01628_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__mux2_1
X_07778_ _00965_ _01574_ _01830_ _01832_ _01569_ VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__a221o_1
X_06729_ _00740_ _00857_ _00535_ VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__a21oi_1
X_09517_ Oset\[1\]\[5\] _03024_ VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_104_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09448_ _03357_ VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09379_ _03288_ _03289_ VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11410_ _05311_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__inv_2
X_12390_ _06131_ net21 VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_50_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11341_ _05241_ _05233_ VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11272_ _05163_ _05168_ _00626_ _02096_ _05173_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__a311o_2
XTAP_TAPCELL_ROW_72_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13011_ clknet_leaf_46_clk _00454_ VGND VGND VPWR VPWR Qset\[3\]\[2\] sky130_fd_sc_hd__dfxtp_2
X_10223_ _04128_ _04129_ VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10154_ Oset\[3\]\[14\] _02787_ _02525_ _04060_ VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__o211a_1
X_10085_ _03991_ _03963_ VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_58_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10987_ _04881_ Qset\[1\]\[12\] _04042_ _04889_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12726_ clknet_leaf_53_clk _00169_ VGND VGND VPWR VPWR H\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12657_ clknet_leaf_26_clk _00107_ VGND VGND VPWR VPWR H\[3\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_11608_ _03770_ _05500_ _05501_ _05507_ _01156_ VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__o221a_1
X_12588_ clknet_leaf_27_clk _00038_ VGND VGND VPWR VPWR Qset\[0\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11539_ _04690_ _04744_ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08750_ _02662_ _02663_ _02539_ VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__nand3_1
X_07701_ result_reg_not\[6\] _01633_ _01759_ VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__a21o_1
X_08681_ _02595_ _00580_ VGND VGND VPWR VPWR _02596_ sky130_fd_sc_hd__nand2_1
X_07632_ _01690_ _01595_ _01692_ _01569_ _01693_ VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__a311o_1
XFILLER_0_88_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07563_ _01623_ _01627_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_75_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09302_ _03209_ _03212_ VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__nand2_1
X_07494_ _01557_ _01558_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__nand2_2
X_06514_ _00625_ _00472_ _00648_ VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__and3b_1
XFILLER_0_63_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09233_ _00587_ R1\[1\] VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__nand2_1
X_06445_ shift.Q VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09164_ _00587_ im_reg\[7\] VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__nand2_1
X_08115_ _01627_ _02055_ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__nor2_4
X_06376_ im_reg\[7\] _00486_ VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09095_ _02992_ _02253_ _03004_ _03005_ VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__o211ai_1
X_08046_ _02036_ VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09997_ _02949_ _03897_ _03899_ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__or3_1
X_08948_ _02653_ _02860_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__nor2_1
X_08879_ _02562_ Qset\[1\]\[2\] VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__nand2_1
X_10910_ _00710_ _04690_ _04813_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__o21ai_2
X_11890_ _05668_ _01602_ VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_55_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10841_ _04308_ _04744_ VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10772_ _04282_ Qset\[1\]\[11\] _03345_ _04675_ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12511_ _06219_ _00490_ VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12442_ _06174_ _06175_ _06138_ VGND VGND VPWR VPWR _06176_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12373_ net24 _06113_ _06117_ net25 _06108_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__a311o_1
XFILLER_0_62_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11324_ _05052_ _05007_ _05224_ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__nand3_1
XFILLER_0_22_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11255_ _05156_ _02473_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__and2_2
X_10206_ _04075_ _04112_ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__nand2_1
X_11186_ _04663_ _04660_ _04693_ VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__o21a_1
X_10137_ _03152_ H\[2\]\[13\] VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10068_ _03049_ _03507_ _03898_ VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__or3_1
XFILLER_0_82_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12709_ clknet_leaf_45_clk _00152_ VGND VGND VPWR VPWR Oset\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09920_ _03826_ _02558_ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09851_ _02556_ VGND VGND VPWR VPWR _03758_ sky130_fd_sc_hd__buf_4
X_06994_ _01111_ VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__clkbuf_1
X_08802_ _02527_ _02182_ _02534_ _02715_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__o211ai_1
X_09782_ _03110_ _03421_ VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08733_ _02647_ VGND VGND VPWR VPWR _02648_ sky130_fd_sc_hd__inv_2
X_08664_ _00004_ VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__buf_6
X_08595_ _02491_ _02510_ VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_52_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07615_ _01677_ VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__clkbuf_1
X_07546_ _01606_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07477_ _00572_ Him VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09216_ _02787_ Qset\[0\]\[5\] _03126_ VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06428_ _00553_ _00562_ VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_60_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06359_ _00497_ _00475_ _00499_ next_PC\[4\] _00478_ VGND VGND VPWR VPWR _00018_
+ sky130_fd_sc_hd__a32o_1
X_09147_ _03057_ _02872_ VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09078_ _02247_ _02161_ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__nand2_1
X_08029_ Oset\[1\]\[8\] _01403_ _02019_ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11040_ _04941_ _04942_ VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__nand2_1
X_12991_ clknet_leaf_6_clk _00434_ VGND VGND VPWR VPWR Qreg2 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11942_ result_reg_Lshift\[5\] _05743_ _05672_ _05787_ VGND VGND VPWR VPWR _00313_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11873_ result_reg_mac\[11\] _05703_ _01149_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10824_ _03866_ VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10755_ _04653_ _04658_ _04654_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__nand3b_1
X_10686_ _04589_ _04590_ VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__nand2_1
X_12425_ _06117_ _06160_ VGND VGND VPWR VPWR _06161_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12356_ _06102_ _00528_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11307_ _04973_ _04924_ VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12287_ _06055_ _00700_ VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11238_ Oset\[1\]\[13\] _04302_ _04303_ VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__o21ai_1
X_11169_ _05070_ _05071_ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07400_ _01276_ _01458_ _01471_ _01472_ VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__a22o_2
XFILLER_0_58_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08380_ _02260_ _02303_ _02250_ _02304_ VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__a211o_1
XFILLER_0_92_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07331_ result_reg_and\[9\] VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07262_ result_reg_add\[5\] _01264_ _01265_ _01341_ VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__o211a_1
X_07193_ _00694_ _01275_ _01276_ VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__a21oi_1
X_09001_ _02912_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09903_ _01538_ _03797_ _03800_ _03809_ VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__a31o_2
X_09834_ _00884_ _02654_ _02753_ _03741_ VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06977_ _01096_ _00735_ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__nand2_1
X_09765_ _03671_ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__inv_2
X_09696_ _03452_ _03599_ _03598_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__o21bai_2
XTAP_TAPCELL_ROW_1_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08716_ Qset\[2\]\[0\] Qset\[3\]\[0\] _00000_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__mux2_1
X_08647_ _02561_ VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_37_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08578_ _02470_ H\[0\]\[14\] VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07529_ _01593_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__clkbuf_4
X_10540_ _00933_ _02654_ _02753_ _04445_ VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__a211o_1
XFILLER_0_36_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10471_ _04376_ VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12210_ _05904_ _05803_ _01243_ _06003_ _05922_ VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12141_ _00525_ _04058_ _05329_ VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_9_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12072_ _02766_ _02769_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__nand2_1
X_11023_ _04925_ VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12974_ clknet_leaf_3_clk _00417_ VGND VGND VPWR VPWR CMD_and sky130_fd_sc_hd__dfxtp_1
X_11925_ _05770_ _05771_ _05710_ _05772_ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__a211o_1
XFILLER_0_87_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11856_ _00811_ _05707_ _05710_ _05717_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__a211o_1
XFILLER_0_74_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11787_ _05669_ VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10807_ _04709_ _04710_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10738_ _02653_ _04642_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12408_ _06132_ _06115_ VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__nand2_1
X_10669_ _04387_ _04386_ VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12339_ _06090_ VGND VGND VPWR VPWR _00407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06900_ _01006_ _00695_ _01022_ _00725_ _00644_ VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__a221o_1
X_07880_ _01691_ result_reg_and\[15\] VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06831_ result_reg_set\[10\] VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__inv_2
X_06762_ result_reg_or\[7\] VGND VGND VPWR VPWR _00890_ sky130_fd_sc_hd__inv_2
X_09550_ _03018_ _02264_ _03458_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09481_ _03386_ _03390_ VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__nor2_1
X_08501_ _02397_ H\[2\]\[11\] VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__nor2_1
X_06693_ shift.left CMD_logic_shift_right _00820_ _00822_ VGND VGND VPWR VPWR _00823_
+ sky130_fd_sc_hd__or4_1
XFILLER_0_53_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08432_ _02354_ net62 _02170_ VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08363_ _02288_ VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__clkbuf_1
X_07314_ _00912_ _00906_ _01174_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__mux2_1
X_08294_ _02218_ _02221_ VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__nand2_2
X_07245_ _00787_ _01266_ _01207_ _01325_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__o211a_1
X_07176_ _01259_ _01255_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09817_ _01537_ _03724_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__nor2_1
X_09748_ _03626_ _03611_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11710_ _01538_ _05597_ _05599_ _05609_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__a31o_2
X_09679_ _03582_ _03587_ _00646_ VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12690_ clknet_leaf_43_clk _00140_ VGND VGND VPWR VPWR Oset\[0\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_11641_ _05535_ _05540_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__xnor2_1
X_11572_ _05471_ _05472_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__nand2_1
Xinput19 instruction_in[11] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_12_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10523_ _04425_ _04426_ _04427_ _04428_ _00647_ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_40_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10454_ _04341_ _04358_ _04359_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10385_ _03760_ Qset\[3\]\[9\] _03761_ _04290_ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_75_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12124_ _04671_ _03866_ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__nand2_1
X_12055_ _02613_ _02615_ _01666_ VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__and3_1
X_11006_ _04907_ _04908_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ clknet_leaf_1_clk _00400_ VGND VGND VPWR VPWR result_reg_set\[12\] sky130_fd_sc_hd__dfxtp_1
X_12888_ clknet_leaf_22_clk _00331_ VGND VGND VPWR VPWR result_reg_Rshift\[7\] sky130_fd_sc_hd__dfxtp_1
X_11908_ result_reg_Lshift\[1\] _05743_ _05672_ _05757_ VGND VGND VPWR VPWR _00309_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11839_ _05705_ VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07030_ _01131_ VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_97_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08981_ _02886_ _02892_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__nand2_1
X_07932_ _01964_ LC\[0\] VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__nand2_1
X_07863_ _01913_ result_reg_mac\[14\] _01540_ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__mux2_1
X_06814_ _00540_ _00933_ _00534_ VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__a21oi_1
X_09602_ _03509_ _03510_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__nand2_1
X_07794_ _01586_ result_reg_sub\[11\] VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__nand2_1
X_09533_ _03439_ VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__inv_2
X_06745_ result_reg_Lshift\[6\] VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__inv_2
X_06676_ _00805_ _00806_ _00643_ VGND VGND VPWR VPWR _00807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09464_ _03366_ _03371_ VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__nand2_1
X_08415_ _02319_ Qset\[2\]\[8\] _02329_ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__o21ai_1
X_09395_ _03304_ _03019_ VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08346_ _02270_ _02147_ _02271_ VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__nand3_1
X_08277_ _02202_ _02203_ _02204_ _02205_ VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__o22a_1
X_07228_ _01309_ _01255_ VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__nand2_1
X_07159_ _01206_ VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10170_ _03136_ Qset\[0\]\[15\] _02526_ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__a21oi_1
X_12811_ clknet_leaf_12_clk _00254_ VGND VGND VPWR VPWR result_reg_add\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_45_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12742_ clknet_leaf_53_clk _00185_ VGND VGND VPWR VPWR H\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12673_ clknet_leaf_28_clk _00123_ VGND VGND VPWR VPWR Oset\[2\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_11624_ _05520_ _05523_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11555_ _05435_ _05455_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__nand2b_1
X_10506_ _04410_ _02092_ _04411_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__nand3_1
X_11486_ _05382_ _05386_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10437_ _04342_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10368_ _04271_ VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__inv_2
X_12107_ _01776_ _05873_ _02115_ _05918_ VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__a211oi_1
X_10299_ _04205_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__inv_2
X_12038_ result_reg_Rshift\[10\] _05848_ _05857_ _05862_ VGND VGND VPWR VPWR _00334_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06530_ _00664_ VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_34_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06461_ _00579_ _00595_ VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__or2b_1
XFILLER_0_34_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08200_ _02127_ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__buf_4
XFILLER_0_28_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06392_ _00526_ VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09180_ _03088_ _03090_ VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__nand2_2
XFILLER_0_16_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08131_ H\[0\]\[7\] _01781_ _02075_ VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08062_ _01781_ H\[2\]\[7\] _02038_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07013_ _01004_ Qset\[1\]\[11\] _01108_ VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08964_ _02561_ Oset\[1\]\[3\] VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__nand2_1
X_07915_ _01953_ VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__clkbuf_1
X_08895_ _02807_ _02552_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__nand2_1
X_07846_ _01894_ _01897_ _01612_ VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__mux2_1
X_07777_ _01571_ _00551_ _01831_ _01667_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__o2bb2a_1
X_06728_ result_reg_add\[6\] VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__inv_2
X_09516_ _03021_ Oset\[0\]\[5\] VGND VGND VPWR VPWR _03426_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09447_ _03355_ _03259_ _03356_ VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_104_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06659_ _00788_ _00789_ _00730_ VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09378_ _03286_ _03282_ _03284_ VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__nand3_1
XFILLER_0_19_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08329_ _02241_ _02253_ _02254_ _02255_ VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_34_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11340_ _05233_ _05241_ VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11271_ _05170_ _05172_ _00626_ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__a21oi_1
X_13010_ clknet_leaf_46_clk _00453_ VGND VGND VPWR VPWR Qset\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10222_ _04127_ _04123_ VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__nand2_1
X_10153_ _02523_ _02483_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_58_Left_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10084_ _03421_ _03876_ VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10986_ _04881_ _02432_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12725_ clknet_leaf_49_clk _00168_ VGND VGND VPWR VPWR H\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_12656_ clknet_leaf_26_clk _00106_ VGND VGND VPWR VPWR H\[3\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_67_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11607_ _02163_ _05506_ VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__nor2_1
X_12587_ clknet_leaf_28_clk _00037_ VGND VGND VPWR VPWR Qset\[0\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11538_ _03233_ _04345_ _05158_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__nor3_1
XFILLER_0_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11469_ _05369_ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_76_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07700_ result_reg_Rshift\[6\] _01672_ _01607_ _01758_ VGND VGND VPWR VPWR _01759_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08680_ _02588_ _02594_ VGND VGND VPWR VPWR _02595_ sky130_fd_sc_hd__nand2_1
X_07631_ result_reg_or\[3\] _01595_ VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07562_ R3\[0\] _01612_ _01625_ _01626_ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__a22o_2
XFILLER_0_75_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06513_ _00647_ _00626_ Qreg3 VGND VGND VPWR VPWR _00648_ sky130_fd_sc_hd__and3_1
X_09301_ _03210_ _03211_ _03207_ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_85_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07493_ _00550_ _00598_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06444_ _00577_ _00578_ VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__nand2_1
X_09232_ _03134_ _03142_ VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06375_ _00511_ _00512_ _00486_ VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__a21bo_1
X_09163_ _03068_ _03073_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08114_ _02073_ VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09094_ _03001_ Oset\[1\]\[4\] VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__nand2_1
X_08045_ _01627_ _01623_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_562 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09996_ _03901_ _03902_ VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__nand2_1
X_08947_ _02858_ _02859_ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__and2_2
X_08878_ _02787_ Qset\[0\]\[2\] VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__nand2_1
X_07829_ _01035_ _01036_ _01544_ VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10840_ _03768_ _04728_ _04743_ _02885_ _00589_ VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__a221oi_4
X_10771_ _03759_ _02409_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12510_ net67 _06220_ _06221_ _06224_ VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12441_ _06147_ _06172_ VGND VGND VPWR VPWR _06175_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12372_ _06115_ _06116_ VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__nand2_2
XFILLER_0_22_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11323_ _05052_ _05007_ _05224_ VGND VGND VPWR VPWR _05225_ sky130_fd_sc_hd__a21o_1
X_11254_ _05150_ _03758_ _00589_ _05155_ VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__a211o_1
X_10205_ _04049_ _02687_ VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11185_ _05086_ _05087_ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__nand2_1
X_10136_ H\[0\]\[13\] H\[1\]\[13\] _02545_ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__mux2_1
X_10067_ _03972_ _03973_ VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10969_ Qset\[1\]\[12\] _04858_ VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12708_ clknet_leaf_3_clk _00012_ VGND VGND VPWR VPWR current_state\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12639_ clknet_leaf_30_clk _00089_ VGND VGND VPWR VPWR Oset\[3\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09850_ _03754_ _03756_ VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__nand2_1
X_06993_ _00722_ Qset\[1\]\[1\] _01109_ VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__mux2_1
X_08801_ _02527_ Oset\[1\]\[1\] VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__nand2_1
X_09781_ _03546_ _03688_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__or2_1
X_08732_ CMD_addition current_state\[6\] VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__nand2_1
X_08663_ _02577_ VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__inv_2
X_08594_ Oset\[0\]\[15\] VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__inv_2
X_07614_ _01676_ H\[3\]\[2\] _01629_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__mux2_1
X_07545_ _01608_ _00659_ _01600_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_52_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07476_ _01540_ VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06427_ _00561_ VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09215_ _02528_ Qset\[1\]\[5\] _02727_ VGND VGND VPWR VPWR _03126_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06358_ _00498_ _00486_ VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__or2_1
X_09146_ _03054_ _03056_ _00581_ VGND VGND VPWR VPWR _03057_ sky130_fd_sc_hd__nand3_1
X_09077_ _02988_ VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__inv_2
X_06289_ _06255_ VGND VGND VPWR VPWR _06256_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08028_ _02027_ VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09979_ _03859_ _02785_ _03050_ VGND VGND VPWR VPWR _03886_ sky130_fd_sc_hd__nand3_2
X_12990_ clknet_leaf_0_clk _00433_ VGND VGND VPWR VPWR shift.Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ _05786_ _05771_ VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _05728_ VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10823_ _04345_ _04495_ VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10754_ _04656_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10685_ _04587_ _04586_ VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__nand2_1
X_12424_ net24 _06266_ _06253_ VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__or3_1
XFILLER_0_23_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12355_ _01146_ VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_17 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11306_ _04994_ _04997_ _04996_ VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12286_ R3\[0\] _06055_ _06044_ _06056_ VGND VGND VPWR VPWR _00388_ sky130_fd_sc_hd__o211a_1
X_11237_ _04832_ Oset\[0\]\[13\] VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__nor2_1
X_11168_ _05069_ _05064_ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__nand2_1
X_10119_ _04025_ _03899_ _04023_ VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11099_ _05000_ _04999_ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07330_ result_reg_not\[9\] _01405_ _01168_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07261_ _01264_ _00841_ VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__nand2_1
X_09000_ _02824_ _02786_ _02911_ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__a21oi_2
X_07192_ _01160_ VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09902_ _03804_ _03808_ _00626_ _00556_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__a31o_1
X_09833_ _02653_ _03740_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06976_ _01092_ _01095_ _00608_ VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__mux2_1
X_09764_ _03669_ _03671_ VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__nand2_1
X_09695_ _03603_ VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08715_ H\[1\]\[0\] _02625_ _00001_ _02629_ VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_1_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _00006_ VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_37_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08577_ H\[1\]\[14\] VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__inv_2
X_07528_ _01567_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07459_ _01527_ _01149_ VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__and2_1
X_10470_ _04374_ _04375_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__nor2_1
X_09129_ Oset\[3\]\[4\] _03025_ _03027_ VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__a21oi_1
X_12140_ _01200_ _04064_ _05324_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__or3_1
XFILLER_0_102_331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12071_ _01578_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11022_ _03233_ _03899_ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12973_ clknet_leaf_3_clk _00416_ VGND VGND VPWR VPWR shift.left sky130_fd_sc_hd__dfxtp_2
X_11924_ result_reg_Lshift\[3\] _05771_ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11855_ _05706_ _03449_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11786_ _00528_ _05668_ VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__nor2_4
XFILLER_0_67_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10806_ _04514_ _04707_ _04511_ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__nand3_1
X_10737_ _04640_ _04641_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_43_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12407_ _06145_ _06146_ _02125_ VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__o21a_1
X_10668_ _04571_ _04572_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__nand2_1
X_10599_ _04503_ _04457_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__nand2_1
X_12338_ _06089_ _01532_ VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12269_ _06032_ _00974_ VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__nand2_1
X_06830_ result_reg_mac\[10\] VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06761_ net14 _00696_ _00888_ VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__o21ai_1
X_06692_ CMD_not _00545_ CMD_and _00821_ VGND VGND VPWR VPWR _00822_ sky130_fd_sc_hd__or4_1
X_09480_ _03389_ VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__inv_2
X_08500_ H\[3\]\[11\] VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__inv_2
X_08431_ _02311_ _02341_ _02140_ _02345_ _02353_ VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__o221ai_4
XTAP_TAPCELL_ROW_34_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08362_ _02287_ net59 _02170_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__mux2_1
X_07313_ result_reg_set\[8\] VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__inv_2
X_08293_ _02219_ _02147_ _02220_ VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__nand3_1
X_07244_ _00788_ _01202_ _01204_ _01324_ VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__a211o_1
XFILLER_0_73_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_12_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07175_ _00700_ _01258_ _01182_ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09816_ _03718_ _03723_ _00647_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06959_ _01074_ _01079_ VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__nand2_1
X_09747_ _03625_ _03627_ _03654_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__nand3_1
XFILLER_0_68_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09678_ _03583_ _03584_ _03026_ _03585_ _03586_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__a32o_1
X_08629_ _02527_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__buf_6
XFILLER_0_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11640_ _05538_ _05539_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__nand2_1
X_11571_ _04955_ _02096_ VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_30_Left_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10522_ Oset\[1\]\[9\] _03792_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10453_ _04357_ _04343_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__nand2_1
X_10384_ _03760_ _02357_ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_75_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12123_ _01831_ _05873_ _02115_ _05931_ VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_20_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12054_ _05872_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11005_ _04906_ _04900_ VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_48_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12956_ clknet_leaf_14_clk _00399_ VGND VGND VPWR VPWR result_reg_set\[11\] sky130_fd_sc_hd__dfxtp_1
X_12887_ clknet_leaf_23_clk _00330_ VGND VGND VPWR VPWR result_reg_Rshift\[6\] sky130_fd_sc_hd__dfxtp_1
X_11907_ _05756_ _05743_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_86_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _02646_ _05703_ _05634_ _05704_ VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__a211o_1
XFILLER_0_74_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11769_ _05627_ _01016_ _02115_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_40_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08980_ _02891_ _02572_ _00586_ VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__a21oi_1
X_07931_ _01963_ _00474_ VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__nand2_4
XFILLER_0_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07862_ _01593_ _01905_ _01912_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__o21ai_1
X_06813_ result_reg_or\[9\] VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09601_ _03508_ _03475_ _03476_ VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__nand3b_1
X_07793_ _01581_ result_reg_add\[11\] VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__nand2_1
X_09532_ _03418_ _02092_ _03419_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__nand3_1
X_06744_ result_reg_not\[6\] VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06675_ result_reg_Lshift\[4\] VGND VGND VPWR VPWR _00806_ sky130_fd_sc_hd__inv_2
X_09463_ _03370_ _03275_ _03372_ VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__nand3_1
X_08414_ Qset\[3\]\[8\] _02260_ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__nor2_1
X_09394_ _03303_ VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08345_ _02141_ Qset\[1\]\[5\] VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_31_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08276_ Oset\[1\]\[2\] _02129_ _02135_ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__o21ai_1
X_07227_ _01306_ _01308_ _01182_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07158_ _01198_ VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07089_ _01173_ VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__buf_4
X_12810_ clknet_leaf_12_clk _00253_ VGND VGND VPWR VPWR result_reg_add\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12741_ clknet_leaf_49_clk _00184_ VGND VGND VPWR VPWR H\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12672_ clknet_leaf_34_clk _00122_ VGND VGND VPWR VPWR Oset\[2\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11623_ _05521_ _05522_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_22_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11554_ _05436_ _05454_ VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10505_ _04345_ _02096_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__nand2_1
X_11485_ _05384_ _05385_ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_40_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10436_ _03899_ _04309_ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10367_ _04266_ _04269_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__nor2_1
X_12106_ _05915_ _05878_ _05916_ _05917_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__and4_1
X_10298_ _03613_ _03350_ _04204_ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__o21ai_1
X_12037_ _05818_ _05851_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12939_ clknet_leaf_22_clk _00382_ VGND VGND VPWR VPWR result_reg_not\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06460_ _00594_ _00528_ _00550_ VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06391_ _00523_ _00525_ VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__nor2_2
XFILLER_0_43_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08130_ _02082_ VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_99_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08061_ _02045_ VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07012_ _01120_ VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08963_ _02874_ _02226_ VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07914_ Oset\[2\]\[10\] _01437_ _01941_ VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__mux2_1
X_08894_ _02801_ _02803_ _02806_ VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__o21ai_4
X_07845_ result_reg_not\[13\] _01600_ _01896_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07776_ result_reg_and\[10\] VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__inv_2
X_06727_ result_reg_mac\[6\] VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__inv_2
X_09515_ H\[1\]\[5\] _03033_ _02840_ _03424_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__a211o_1
XFILLER_0_91_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09446_ _03252_ _03250_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_104_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06658_ result_reg_add\[4\] VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09377_ _03285_ _03287_ VGND VGND VPWR VPWR _03288_ sky130_fd_sc_hd__nand2_1
X_06589_ _00722_ Qset\[0\]\[1\] _00687_ VGND VGND VPWR VPWR _00723_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08328_ _02241_ Oset\[1\]\[4\] VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_104_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08259_ H\[0\]\[1\] VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11270_ _02469_ _04855_ _05171_ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_72_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10221_ _04123_ _04127_ VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__or2_1
X_10152_ _02162_ _04058_ _02796_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__o21ai_1
X_10083_ _03965_ _03989_ VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_58_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12724_ clknet_leaf_30_clk _00167_ VGND VGND VPWR VPWR Oset\[1\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10985_ Qset\[2\]\[12\] Qset\[3\]\[12\] _04729_ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12655_ clknet_leaf_33_clk _00105_ VGND VGND VPWR VPWR H\[3\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_11606_ _05502_ _05503_ _04303_ _05504_ _05505_ VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__a32o_1
XFILLER_0_65_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12586_ clknet_leaf_29_clk _00036_ VGND VGND VPWR VPWR Qset\[0\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11537_ _05182_ _05180_ _05179_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11468_ _05362_ _05368_ VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11399_ _05300_ _02160_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__nand2_1
X_10419_ _04260_ _04324_ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_2_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07630_ _01691_ result_reg_and\[3\] VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__nand2_1
X_07561_ _00498_ _01541_ _01606_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__o21a_1
X_06512_ _00646_ VGND VGND VPWR VPWR _00647_ sky130_fd_sc_hd__clkbuf_8
X_09300_ _03201_ _03199_ VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__nand2_1
X_07492_ _00557_ _01556_ VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06443_ CMD_not VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09231_ _03141_ _02573_ _00587_ VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__a21oi_1
X_06374_ next_PC\[7\] _00508_ VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__or2_1
X_09162_ _03072_ _02572_ _00586_ VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08113_ _01938_ H\[1\]\[15\] _02056_ VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09093_ _02591_ VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__buf_6
XFILLER_0_31_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08044_ _02035_ VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09995_ _03900_ _03894_ _03895_ VGND VGND VPWR VPWR _03902_ sky130_fd_sc_hd__nand3b_1
X_08946_ _02857_ _02855_ _02856_ VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__nand3_1
X_08877_ _02788_ _02525_ _02789_ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__nand3_2
X_07828_ _01880_ VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_55_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07759_ _01808_ _01541_ _01814_ _01612_ VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10770_ _04282_ Qset\[3\]\[11\] _03761_ _04673_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09429_ _03337_ _03338_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__nand2_1
X_12440_ _06104_ _06140_ VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12371_ net20 net21 VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__nor2_2
XFILLER_0_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11322_ _05222_ _05223_ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__nand2_1
X_11253_ _03758_ _05154_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__nor2_1
X_10204_ _03115_ _04110_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11184_ _05085_ _05061_ VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10135_ _02560_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__buf_4
XFILLER_0_89_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10066_ _03971_ _03970_ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__nand2_1
X_10968_ _04856_ Qset\[0\]\[12\] _04862_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__a21oi_1
X_12707_ clknet_leaf_2_clk _00011_ VGND VGND VPWR VPWR current_state\[5\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_57_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12638_ clknet_leaf_30_clk _00088_ VGND VGND VPWR VPWR Oset\[3\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10899_ Qset\[3\]\[11\] _03792_ _03795_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12569_ clknet_leaf_38_clk _00019_ VGND VGND VPWR VPWR next_PC\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08800_ _02161_ _02711_ _02713_ VGND VGND VPWR VPWR _02714_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09780_ _03076_ _03421_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__nand2_1
X_06992_ _01110_ VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__clkbuf_1
X_08731_ _02645_ VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08662_ _02575_ _02576_ VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__nand2_2
X_07613_ _01671_ _01675_ _01613_ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__mux2_4
XFILLER_0_72_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08593_ _02491_ Oset\[3\]\[15\] _02374_ _02508_ VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__a211o_1
X_07544_ result_reg_Rshift\[0\] _01608_ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_52_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07475_ _00625_ _01539_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__nor2_4
XFILLER_0_91_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06426_ _00560_ VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__clkbuf_4
X_09214_ _02523_ Qset\[2\]\[5\] _03124_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06357_ R1\[0\] VGND VGND VPWR VPWR _00498_ sky130_fd_sc_hd__clkbuf_8
X_09145_ _02528_ Qset\[1\]\[7\] _02727_ _03055_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__a211o_1
X_09076_ _00762_ _02654_ _02753_ _02987_ VGND VGND VPWR VPWR _02988_ sky130_fd_sc_hd__a211o_1
X_06288_ net20 net21 VGND VGND VPWR VPWR _06255_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08027_ Oset\[1\]\[7\] _01385_ _02019_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09978_ _03883_ _03884_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__nand2_1
X_08929_ H\[1\]\[2\] _02836_ _02840_ _02841_ VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__a211o_1
X_11940_ _05769_ _05785_ _05755_ VGND VGND VPWR VPWR _05786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ _00955_ _05707_ _05710_ _05727_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10822_ _04558_ _04539_ _04557_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_80_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10753_ _04653_ _04655_ _04656_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10684_ _04588_ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__inv_2
X_12423_ _06126_ _06158_ _04827_ _06159_ VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12354_ _06097_ CMD_addition _06066_ _06101_ VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11305_ _05205_ _05206_ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12285_ _06055_ _01170_ VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11236_ Oset\[3\]\[13\] _04302_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__nor2_1
X_11167_ _05064_ _05069_ VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10118_ _03789_ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__inv_2
X_11098_ _04999_ _05000_ VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10049_ _03951_ _03955_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__nor2_2
XFILLER_0_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07260_ _01338_ _01187_ _01192_ _01339_ VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__a211o_1
X_07191_ _01220_ VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09901_ _03805_ _03794_ _00621_ _03807_ VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__a211o_1
XFILLER_0_41_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09832_ _03738_ _03739_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__and2_2
X_09763_ _03670_ _03228_ VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__nand2_1
X_06975_ _01086_ _01094_ _00613_ VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__mux2_1
X_08714_ _02625_ _02155_ VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__nor2_1
X_09694_ _00857_ _02654_ _02753_ _03602_ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_1_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08645_ _02525_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_65_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08576_ _02490_ _02491_ _02374_ _02492_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__a211o_1
X_07527_ _01209_ _01577_ _01591_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_91_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_558 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07458_ R2\[0\] net27 current_state\[2\] VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06409_ result_reg_sub\[0\] _00540_ VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__or2_1
X_07389_ _01010_ _01266_ _01299_ _01461_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09128_ Oset\[1\]\[4\] _03033_ VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_9_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09059_ Qset\[1\]\[3\] _02836_ VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__nand2_1
X_12070_ _00715_ _05873_ _05775_ _05887_ VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__a211oi_1
X_11021_ _04854_ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_99_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12972_ clknet_leaf_7_clk _00415_ VGND VGND VPWR VPWR CMD_logic_shift_right sky130_fd_sc_hd__dfxtp_2
X_11923_ _05741_ VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__clkbuf_4
X_11854_ _05716_ VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__inv_2
X_10805_ _04647_ _04708_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__nand2_1
X_11785_ _05667_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10736_ _04639_ _04638_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10667_ _04532_ _04534_ _04569_ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__nand3_1
X_12406_ _06140_ _06138_ _06112_ _01146_ VGND VGND VPWR VPWR _06146_ sky130_fd_sc_hd__and4_1
XFILLER_0_23_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10598_ _04497_ _04501_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__nand2_1
X_12337_ im_reg\[6\] net31 _01146_ VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12268_ _06039_ _05805_ _06044_ _06045_ VGND VGND VPWR VPWR _00381_ sky130_fd_sc_hd__o211a_1
X_11219_ _04824_ _04639_ _04638_ VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__nand3_1
X_12199_ _05937_ _05993_ _05994_ _05904_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06760_ _00887_ _00735_ VGND VGND VPWR VPWR _00888_ sky130_fd_sc_hd__nand2_1
X_06691_ CMD_set _00697_ _00593_ VGND VGND VPWR VPWR _00821_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_62_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08430_ _02349_ _02352_ _01553_ VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_34_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08361_ _02126_ _02273_ _02140_ _02280_ _02286_ VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__o221ai_2
X_07312_ net15 _01255_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08292_ _02131_ Qset\[1\]\[3\] VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__nand2_1
X_07243_ result_reg_add\[4\] _01202_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07174_ _00701_ _01257_ _01177_ VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09815_ _03719_ _03720_ _03027_ _03721_ _03722_ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__a32o_1
XFILLER_0_94_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06958_ _01075_ _00654_ _00656_ _01078_ _00665_ VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__a221o_1
X_09746_ _03653_ VGND VGND VPWR VPWR _03654_ sky130_fd_sc_hd__inv_2
X_09677_ _03021_ Qset\[2\]\[6\] VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__nand2_1
X_06889_ result_reg_and\[12\] _00561_ _00552_ VGND VGND VPWR VPWR _01012_ sky130_fd_sc_hd__o21ai_1
X_08628_ _02161_ _02538_ _02542_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__o21ai_1
X_08559_ Qset\[2\]\[14\] VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11570_ _05470_ _04830_ VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10521_ _04414_ Oset\[0\]\[9\] _03798_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10452_ _04343_ _04357_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__or2_1
X_10383_ _02363_ _02163_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_75_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12122_ _05927_ _05929_ _05930_ _05871_ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__and4_1
X_12053_ _05871_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__inv_2
X_11004_ _04900_ _04906_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__or2_1
X_12955_ clknet_leaf_15_clk _00398_ VGND VGND VPWR VPWR result_reg_set\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_48_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11906_ _05748_ _05753_ _05755_ VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12886_ clknet_leaf_23_clk _00329_ VGND VGND VPWR VPWR result_reg_Rshift\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ result_reg_mac\[0\] _05702_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11768_ _05626_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10719_ Oset\[3\]\[10\] _03791_ _03027_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__a21oi_1
X_11699_ H\[1\]\[15\] _04858_ _04862_ _05598_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_11_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07930_ _06284_ _01962_ VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07861_ _01909_ _01572_ _01910_ _01568_ _01911_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__a311o_1
XFILLER_0_47_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06812_ net16 _00696_ _00937_ VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__o21ai_1
X_07792_ _01843_ _01658_ _01844_ _01845_ VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__a31o_1
X_09600_ _03477_ _03508_ VGND VGND VPWR VPWR _03509_ sky130_fd_sc_hd__nand2_1
X_06743_ _00856_ _00695_ _00871_ _00725_ _00644_ VGND VGND VPWR VPWR _00872_ sky130_fd_sc_hd__a221o_1
X_09531_ _03413_ _00536_ _03414_ VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__nand3_1
XFILLER_0_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06674_ result_reg_Rshift\[4\] VGND VGND VPWR VPWR _00805_ sky130_fd_sc_hd__inv_2
X_09462_ _03362_ _03365_ _03371_ VGND VGND VPWR VPWR _03372_ sky130_fd_sc_hd__nand3_1
XFILLER_0_93_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08413_ _02336_ VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__clkbuf_1
X_09393_ _02734_ _03079_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__nand2_1
X_08344_ _02230_ Qset\[0\]\[5\] VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08275_ _02131_ Oset\[0\]\[2\] VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07226_ _00765_ _01307_ _01177_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07157_ _01227_ _01241_ _00669_ _01159_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_14_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07088_ _00538_ _01172_ VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__nand2_4
X_09729_ _03001_ Qset\[0\]\[7\] VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_45_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12740_ clknet_leaf_26_clk _00183_ VGND VGND VPWR VPWR H\[2\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_12671_ clknet_leaf_38_clk _00121_ VGND VGND VPWR VPWR Oset\[2\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_11622_ _04073_ _05158_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11553_ _05452_ _05453_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__nand2_1
X_10504_ _04408_ _04409_ _00710_ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__nand3_1
X_11484_ _05383_ _05259_ VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__nand2_1
X_10435_ _04024_ _04021_ VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12105_ _00525_ _03639_ _05789_ VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__or3_1
X_10366_ _04266_ _04269_ _04271_ VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__o21ai_1
X_10297_ _03505_ _03462_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__nand2_1
X_12036_ result_reg_Rshift\[9\] _05848_ _05857_ _05861_ VGND VGND VPWR VPWR _00333_
+ sky130_fd_sc_hd__o211a_1
X_12938_ clknet_leaf_22_clk _00381_ VGND VGND VPWR VPWR result_reg_not\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12869_ clknet_leaf_19_clk _00312_ VGND VGND VPWR VPWR result_reg_Lshift\[4\] sky130_fd_sc_hd__dfxtp_1
X_06390_ _00524_ VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_55_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08060_ _01761_ H\[2\]\[6\] _02038_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07011_ _00979_ Qset\[1\]\[10\] _01108_ VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08962_ _00006_ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__clkbuf_4
X_07913_ _01952_ VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__clkbuf_1
X_08893_ _02804_ _02525_ _02805_ VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__nand3_1
X_07844_ result_reg_Rshift\[13\] _01672_ _01601_ _01895_ VGND VGND VPWR VPWR _01896_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07775_ _01827_ _01663_ _01828_ _01829_ VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__a31o_1
X_06726_ _00855_ VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__clkbuf_1
X_09514_ _03033_ _02281_ VGND VGND VPWR VPWR _03424_ sky130_fd_sc_hd__nor2_1
X_06657_ result_reg_sub\[4\] VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09445_ _03250_ _03252_ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06588_ _00645_ _00693_ _00721_ VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__o21ai_4
X_09376_ _03286_ VGND VGND VPWR VPWR _03287_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08327_ _02147_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08258_ _02129_ _02186_ _02135_ _02187_ VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__a211o_1
X_07209_ _01290_ _01193_ _01191_ _01291_ VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__a211o_1
X_08189_ _02119_ _02120_ VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10220_ _04115_ _04124_ _04126_ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10151_ _04055_ _04057_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__nand2_2
X_10082_ _03349_ _03868_ VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_58_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10984_ _03770_ _04886_ _01156_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_83_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12723_ clknet_leaf_30_clk _00166_ VGND VGND VPWR VPWR Oset\[1\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12654_ clknet_leaf_33_clk _00104_ VGND VGND VPWR VPWR H\[3\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_11605_ Qset\[3\]\[15\] _04302_ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__or2_1
X_12585_ clknet_leaf_35_clk _00035_ VGND VGND VPWR VPWR Qset\[0\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11536_ _04926_ _05379_ VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11467_ _05363_ _05367_ VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11398_ _00820_ _04974_ _05299_ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10418_ _04322_ _04323_ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__nand2_1
X_10349_ _04254_ _04255_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__and2_2
X_12019_ _05847_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07560_ R0\[0\] _01568_ _01540_ _01624_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06511_ Oreg3 VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__inv_2
X_07491_ _01555_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09230_ _03135_ _03137_ _03138_ _03140_ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__a31o_2
X_06442_ _00545_ _00576_ VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06373_ _00508_ next_PC\[7\] VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09161_ _03069_ _03070_ _03071_ _02526_ VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__a22oi_4
X_08112_ _02072_ VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__clkbuf_1
X_09092_ _03001_ _02249_ _02991_ _03002_ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__o211ai_1
X_08043_ Oset\[1\]\[15\] _01525_ _02018_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09994_ _03896_ _03900_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08945_ _02855_ _02856_ _02857_ VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08876_ _02562_ Qset\[3\]\[2\] VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07827_ _01879_ H\[3\]\[12\] _01628_ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__mux2_1
X_07758_ _01811_ _01746_ _01812_ _01593_ _01813_ VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_55_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06709_ _00838_ VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07689_ _01744_ _01635_ _01745_ _01747_ VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__a31o_1
XFILLER_0_66_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09428_ _02280_ _00583_ VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09359_ _02828_ _02955_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__nor2_1
X_12370_ net23 _06114_ VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11321_ _05221_ _05220_ VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11252_ _05151_ _05152_ _05153_ _04835_ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__a22o_1
X_11183_ _05061_ _05085_ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__or2_1
X_10203_ _04109_ VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__inv_2
X_10134_ _04031_ _04040_ VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__nand2_1
X_10065_ _03970_ _03971_ VGND VGND VPWR VPWR _03972_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10967_ _04856_ Qset\[2\]\[12\] VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__nand2_1
X_12706_ clknet_leaf_3_clk _00010_ VGND VGND VPWR VPWR current_state\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10898_ Qset\[1\]\[11\] _03792_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__nand2_1
X_12637_ clknet_leaf_28_clk _00087_ VGND VGND VPWR VPWR Oset\[3\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12568_ clknet_leaf_38_clk _00018_ VGND VGND VPWR VPWR next_PC\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12499_ current_state\[1\] _06271_ _06269_ _00631_ VGND VGND VPWR VPWR _06216_ sky130_fd_sc_hd__and4b_1
X_11519_ _05415_ _05419_ VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__xnor2_1
X_06991_ _00668_ Qset\[1\]\[0\] _01109_ VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__mux2_1
X_08730_ _02623_ _02644_ VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__xor2_4
X_08661_ R3\[0\] _00587_ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__nand2_1
X_07612_ result_reg_not\[2\] _01633_ _01674_ VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08592_ _02491_ _02507_ VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__nor2_1
X_07543_ _01603_ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_3_5__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07474_ _00472_ _01538_ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06425_ _00559_ _00526_ VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09213_ _02528_ Qset\[3\]\[5\] _02534_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09144_ _02561_ _02315_ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_32_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06356_ _00495_ _00496_ _00486_ VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__a21bo_1
X_09075_ _02653_ _02986_ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__nor2_1
X_06287_ net23 net24 VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08026_ _02026_ VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09977_ _03882_ _03860_ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__nand2_1
X_08928_ _02688_ _02210_ VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08859_ _02771_ VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__inv_2
X_11870_ _05706_ _04642_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10821_ _03899_ _04691_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10752_ _04494_ _04270_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12422_ _06126_ _00576_ VGND VGND VPWR VPWR _06159_ sky130_fd_sc_hd__nand2_1
X_10683_ _04586_ _04587_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12353_ _06098_ _06099_ _06100_ _06267_ VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12284_ _06054_ VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__buf_2
X_11304_ _05202_ _04947_ _04952_ VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__nand3_1
XFILLER_0_50_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11235_ _04832_ Oset\[2\]\[13\] VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_91_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11166_ _05066_ _05068_ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__nand2_1
X_11097_ _04958_ _04983_ _04986_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__o21a_1
X_10117_ _04023_ _03790_ _03835_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__nand3b_1
X_10048_ _03953_ _03954_ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11999_ _04078_ _04080_ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07190_ _01254_ _01256_ _01260_ _01273_ VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__a31o_1
X_09900_ Qset\[3\]\[8\] _03023_ _03798_ _03806_ VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09831_ _03737_ _03604_ VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06974_ _01093_ _01083_ _00611_ VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__mux2_1
X_09762_ _03218_ _03219_ _03227_ VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__a21o_1
X_08713_ H\[3\]\[0\] _02625_ _02626_ _02627_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__a211o_1
X_09693_ _02653_ _03601_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08644_ _00584_ _02554_ _02558_ VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_1_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ _02491_ H\[2\]\[14\] VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__nor2_1
X_07526_ _01582_ _01585_ _01587_ _01590_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07457_ _01526_ VGND VGND VPWR VPWR _00089_ sky130_fd_sc_hd__clkbuf_1
X_06408_ _00541_ _00542_ _00535_ VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__a21oi_1
X_07388_ _01016_ _01267_ _01263_ _01460_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06339_ _00481_ _00482_ _06285_ VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__o21ai_1
X_09127_ _03022_ Oset\[0\]\[4\] VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__nand2_1
X_09058_ _02632_ Qset\[0\]\[3\] _02840_ VGND VGND VPWR VPWR _02970_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08009_ Oset\[0\]\[15\] _01525_ _02000_ VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11020_ _03899_ _04691_ _04753_ _04751_ VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__o31a_1
X_12971_ clknet_leaf_1_clk _00414_ VGND VGND VPWR VPWR CMD_mul_accumulation sky130_fd_sc_hd__dfxtp_1
X_11922_ _05755_ _05753_ _05765_ _05769_ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__o22a_1
X_11853_ _00785_ _05707_ _05710_ _05715_ VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10804_ _04707_ VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11784_ _06269_ _05666_ VGND VGND VPWR VPWR _05667_ sky130_fd_sc_hd__nor2_2
X_10735_ _04638_ _04639_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__or2_1
X_10666_ _04535_ _04570_ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__nand2_2
XFILLER_0_82_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12405_ _06102_ _00578_ VGND VGND VPWR VPWR _06145_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10597_ _04457_ _04497_ _04501_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__nand3b_2
X_12336_ _06088_ VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__clkbuf_1
X_12267_ _06033_ _00948_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11218_ _05120_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__inv_2
X_12198_ _03647_ _03072_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__nand2_1
X_11149_ _05050_ _05009_ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06690_ _00710_ VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__buf_6
XFILLER_0_53_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08360_ _02283_ _02285_ _01552_ VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_34_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07311_ result_reg_not\[8\] _01387_ _01167_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08291_ _02151_ Qset\[0\]\[3\] VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__nand2_1
X_07242_ result_reg_and\[4\] VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07173_ _00702_ _00703_ _01174_ VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09814_ _03022_ Qset\[2\]\[7\] VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__nand2_1
X_06957_ result_reg_Rshift\[14\] _00753_ _01077_ VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__o21ai_1
X_09745_ _03652_ _03257_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__nand2_1
X_06888_ _01010_ _00745_ VGND VGND VPWR VPWR _01011_ sky130_fd_sc_hd__or2_1
X_09676_ Qset\[3\]\[6\] _03024_ _03026_ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__a21oi_1
X_08627_ _02541_ VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08558_ _02475_ VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__clkbuf_1
X_07509_ _01573_ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08489_ Qset\[0\]\[11\] VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__inv_2
X_10520_ _04414_ Oset\[2\]\[9\] VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10451_ _04355_ _04356_ VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__nand2_1
X_10382_ _04285_ _04287_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__nand2_2
XFILLER_0_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12121_ _00525_ _04552_ _04477_ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__or3_1
XFILLER_0_102_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12052_ _05870_ _00555_ _05667_ VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__and3_2
X_11003_ _04904_ _04905_ VGND VGND VPWR VPWR _04906_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12954_ clknet_leaf_15_clk _00397_ VGND VGND VPWR VPWR result_reg_set\[9\] sky130_fd_sc_hd__dfxtp_1
X_11905_ _05754_ VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__clkbuf_4
X_12885_ clknet_leaf_19_clk _00328_ VGND VGND VPWR VPWR result_reg_Rshift\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_86_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _05702_ VGND VGND VPWR VPWR _05703_ sky130_fd_sc_hd__buf_4
XFILLER_0_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11767_ _05654_ VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10718_ Oset\[1\]\[10\] _03791_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11698_ _04858_ _02514_ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10649_ _04547_ _04553_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_11_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12319_ _01447_ _06058_ VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07860_ result_reg_or\[14\] _01595_ VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__nor2_1
X_06811_ _00936_ _00735_ VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__nand2_1
X_07791_ net3 _01746_ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06742_ _00739_ _00863_ _00864_ _00869_ _00870_ VGND VGND VPWR VPWR _00871_ sky130_fd_sc_hd__a32o_1
X_09530_ _03415_ _03420_ _03439_ VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09461_ _03369_ VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__inv_2
X_06673_ result_reg_not\[4\] VGND VGND VPWR VPWR _00804_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08412_ _02335_ net61 _02170_ VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__mux2_1
X_09392_ _03301_ _03240_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08343_ _02267_ _02143_ _02268_ VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__nand3_1
X_08274_ _02127_ Oset\[2\]\[2\] _00003_ VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07225_ _00770_ _00762_ _01174_ VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07156_ _01239_ _01214_ _01240_ _01159_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__a31o_1
X_07087_ _01171_ VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07989_ Oset\[0\]\[5\] _01349_ _02001_ VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__mux2_1
X_09728_ _02992_ Qset\[2\]\[7\] _02991_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09659_ _03566_ _02092_ _03567_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__nand3_1
X_12670_ clknet_leaf_37_clk _00120_ VGND VGND VPWR VPWR Oset\[2\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_11621_ _04095_ _04924_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11552_ _05451_ _05437_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11483_ _05259_ _05383_ VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__nor2_1
X_10503_ _04335_ _03746_ _04336_ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__nand3_1
X_10434_ _04040_ _04028_ VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__nand2_1
X_10365_ _03789_ _04270_ VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__nand2_1
X_12104_ _01200_ _03063_ _03632_ VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__or3_1
X_10296_ _03612_ _04202_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__nor2_1
X_12035_ _05814_ _05851_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12937_ clknet_leaf_22_clk _00380_ VGND VGND VPWR VPWR result_reg_not\[8\] sky130_fd_sc_hd__dfxtp_1
X_12868_ clknet_leaf_23_clk _00311_ VGND VGND VPWR VPWR result_reg_Lshift\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11819_ _04527_ _04605_ _05677_ _05691_ VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12799_ clknet_leaf_40_clk _00242_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_99_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07010_ _01119_ VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08961_ _02870_ _02872_ VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__nand2_1
X_07912_ Oset\[2\]\[9\] _01420_ _01942_ VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__mux2_1
X_08892_ _02798_ Oset\[3\]\[2\] VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__nand2_1
X_07843_ _01716_ _01050_ VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__nand2_1
X_07774_ result_reg_mul\[10\] _01688_ _01589_ VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09513_ H\[2\]\[5\] _03022_ _03422_ VGND VGND VPWR VPWR _03423_ sky130_fd_sc_hd__a21o_1
X_06725_ _00854_ Qset\[0\]\[5\] _00687_ VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__mux2_1
X_06656_ result_reg_mul\[4\] VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__inv_2
X_09444_ _03352_ _03353_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06587_ _00694_ _00695_ _00720_ _00628_ _00644_ VGND VGND VPWR VPWR _00721_ sky130_fd_sc_hd__a221o_1
X_09375_ _02985_ _02982_ _03233_ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08326_ Oset\[0\]\[4\] VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08257_ H\[3\]\[1\] _02129_ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07208_ net9 _01186_ VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__nor2_1
X_08188_ CMD_not CMD_logic_shift_right VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07139_ _00498_ _01220_ _01159_ _01223_ VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_18_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10150_ _02565_ _02476_ _04056_ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10081_ _03858_ _03506_ _03050_ VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_58_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10983_ _04882_ _04883_ _04884_ _04885_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_27_Left_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12722_ clknet_leaf_28_clk _00165_ VGND VGND VPWR VPWR Oset\[1\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_83_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12653_ clknet_leaf_40_clk _00103_ VGND VGND VPWR VPWR H\[3\]\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_37_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11604_ _05335_ Qset\[2\]\[15\] _04835_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__o21a_1
X_12584_ clknet_leaf_33_clk _00034_ VGND VGND VPWR VPWR Qset\[0\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11535_ _05185_ _05176_ _05184_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_36_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11466_ _05365_ _05366_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__nor2b_1
XTAP_TAPCELL_ROW_94_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11397_ _05229_ _05298_ _00820_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__nand3_1
X_10417_ _04318_ _03411_ _04319_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10348_ _03812_ _03814_ _04253_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__nand3_1
X_10279_ _04185_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__inv_2
X_12018_ result_reg_Rshift\[2\] _05848_ _05808_ _05850_ VGND VGND VPWR VPWR _00326_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Left_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06510_ _00644_ VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__inv_2
X_07490_ _01554_ _00531_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06441_ CMD_set VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09160_ H\[2\]\[7\] H\[3\]\[7\] _02561_ VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06372_ _00505_ _00475_ _00510_ next_PC\[6\] _00478_ VGND VGND VPWR VPWR _00020_
+ sky130_fd_sc_hd__a32o_1
X_08111_ _01918_ H\[1\]\[14\] _02056_ VGND VGND VPWR VPWR _02072_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_54_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09091_ _03001_ Oset\[3\]\[4\] VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08042_ _02034_ VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09993_ _03897_ _03205_ _03899_ VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__or3_1
XFILLER_0_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08944_ _02749_ _02744_ VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__nand2_1
X_08875_ _02787_ Qset\[2\]\[2\] VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__nand2_1
X_07826_ _01875_ _01878_ _01612_ VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__mux2_1
X_07757_ net16 _01746_ VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06708_ _00837_ _00730_ _00607_ VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_55_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07688_ net13 _01746_ VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__nor2_1
X_06639_ _00770_ _00762_ _00730_ VGND VGND VPWR VPWR _00771_ sky130_fd_sc_hd__mux2_1
X_09427_ _03331_ _01155_ _03336_ VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__nand3_1
XFILLER_0_81_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09358_ _03264_ _03268_ VGND VGND VPWR VPWR _03269_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08309_ _02233_ _02236_ _01551_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11320_ _05220_ _05221_ VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09289_ _03199_ VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11251_ H\[2\]\[13\] H\[3\]\[13\] _04832_ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__mux2_1
X_10202_ _03758_ _04108_ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__nor2_2
X_11182_ _05083_ _05084_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__and2_1
X_10133_ _04038_ _04039_ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__nand2_2
X_10064_ _03933_ _03929_ VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10966_ Qset\[3\]\[12\] _04858_ _04859_ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12705_ clknet_leaf_5_clk _00013_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dfxtp_1
X_10897_ _04414_ Qset\[0\]\[11\] VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__nand2_1
X_12636_ clknet_leaf_34_clk _00086_ VGND VGND VPWR VPWR Oset\[3\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12567_ clknet_leaf_38_clk _00017_ VGND VGND VPWR VPWR next_PC\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11518_ _05417_ _05418_ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__and2b_1
X_12498_ _06215_ VGND VGND VPWR VPWR _00441_ sky130_fd_sc_hd__clkbuf_1
X_11449_ Oset\[3\]\[14\] _04857_ _04859_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06990_ _01108_ VGND VGND VPWR VPWR _01109_ sky130_fd_sc_hd__clkbuf_8
X_08660_ _02559_ _02574_ VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__nand2_1
X_07611_ result_reg_Rshift\[2\] _01672_ _01607_ _01673_ VGND VGND VPWR VPWR _01674_
+ sky130_fd_sc_hd__o211a_1
X_08591_ Oset\[2\]\[15\] VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07542_ _01601_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07473_ _01537_ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__buf_4
X_06424_ _00472_ _00555_ _00556_ _00558_ VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__and4_2
XFILLER_0_63_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09212_ _03122_ _02552_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09143_ _02528_ Qset\[3\]\[7\] _02534_ _03053_ VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__a211o_1
X_06355_ next_PC\[4\] _00491_ VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06286_ net25 VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__inv_2
X_09074_ _02984_ _02985_ VGND VGND VPWR VPWR _02986_ sky130_fd_sc_hd__and2_2
XFILLER_0_44_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08025_ Oset\[1\]\[6\] _01368_ _02019_ VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09976_ _03860_ _03882_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__or2_1
X_08927_ _00001_ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__buf_4
X_08858_ _02770_ _01153_ VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__nand2_1
X_07809_ result_reg_mul\[12\] _01679_ _01656_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_68_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08789_ _01536_ _02690_ _02692_ _00548_ _02702_ VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__a311o_1
XFILLER_0_79_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10820_ _04571_ _04568_ VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10751_ _04654_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12421_ _06154_ _06122_ _06157_ VGND VGND VPWR VPWR _06158_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10682_ _04376_ _04373_ _04381_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__o21a_1
X_12352_ net23 VGND VGND VPWR VPWR _06100_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12283_ _06052_ _06053_ VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__nand2_2
X_11303_ _05203_ _05204_ VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11234_ _05136_ VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_78_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11165_ _05067_ _03688_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__nand2_1
X_11096_ _04994_ _04998_ VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__xnor2_1
X_10116_ _04021_ _04022_ VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__nand2_1
X_10047_ _03904_ _03917_ _03913_ VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__nand3b_1
X_11998_ result_reg_Lshift\[13\] _05743_ _05808_ _05835_ VGND VGND VPWR VPWR _00321_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10949_ _03768_ _04836_ _04850_ _04851_ VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12619_ clknet_leaf_28_clk _00069_ VGND VGND VPWR VPWR Qset\[2\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09830_ _03604_ _03737_ VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06973_ result_reg_sub\[15\] VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__inv_2
X_09761_ _03667_ _03668_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__nand2_1
X_08712_ _02625_ _02152_ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__nor2_1
X_09692_ _03452_ _03600_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__xor2_4
XTAP_TAPCELL_ROW_65_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08643_ _02557_ VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_1_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08574_ _02470_ VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__buf_4
X_07525_ result_reg_mul\[0\] _01585_ _01589_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07456_ Oset\[3\]\[15\] _01525_ _01249_ VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06407_ result_reg_add\[0\] VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__inv_2
X_07387_ result_reg_add\[12\] _01267_ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06338_ next_PC\[1\] next_PC\[0\] VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__nor2_1
X_09126_ _03032_ _03034_ _03027_ _03035_ _03036_ VGND VGND VPWR VPWR _03037_ sky130_fd_sc_hd__a32o_1
XFILLER_0_32_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09057_ _02632_ Qset\[2\]\[3\] VGND VGND VPWR VPWR _02969_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08008_ _02016_ VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09959_ _03862_ _03863_ _02800_ _03864_ _03865_ VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__a32o_2
XFILLER_0_99_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12970_ clknet_leaf_3_clk _00413_ VGND VGND VPWR VPWR Add.sub sky130_fd_sc_hd__dfxtp_1
X_11921_ _05745_ _03169_ _03155_ _05766_ _05768_ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__a221o_2
X_11852_ _05706_ _03293_ VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__nor2_1
X_10803_ _04702_ _04706_ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__nand2_1
X_11783_ _02093_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_52_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10734_ _04255_ _04440_ _04438_ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10665_ _04569_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__inv_2
X_12404_ _06097_ _00545_ _04827_ _06144_ VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10596_ _04498_ _04499_ _04500_ VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__nand3_1
X_12335_ _01534_ _01532_ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__and2_1
X_12266_ _01148_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__clkbuf_4
X_11217_ _05118_ _05119_ VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__nand2_1
X_12197_ _03063_ _03632_ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__nand2_1
Xoutput70 net70 VGND VGND VPWR VPWR instruction_address[5] sky130_fd_sc_hd__clkbuf_1
X_11148_ _05009_ _05050_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__or2_1
X_11079_ _04981_ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07310_ result_reg_Lshift\[8\] result_reg_Rshift\[8\] _01164_ VGND VGND VPWR VPWR
+ _01387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_43_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08290_ _02216_ _02143_ _02217_ VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__nand3_1
X_07241_ _01320_ _01187_ _01192_ _01321_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_14_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07172_ net8 _01255_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_446 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09813_ Qset\[3\]\[7\] _03033_ _03026_ VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__a21oi_1
X_06956_ _00754_ _01076_ VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__nand2_1
X_09744_ _03651_ VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__buf_6
X_06887_ result_reg_mul\[12\] VGND VGND VPWR VPWR _01010_ sky130_fd_sc_hd__inv_2
X_09675_ Qset\[1\]\[6\] _03024_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08626_ _01959_ _00580_ _02540_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_34_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_8
X_08557_ _02474_ net52 _02169_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07508_ _01572_ VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08488_ _02328_ Qset\[3\]\[11\] _02347_ _02407_ VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__a211o_1
X_07439_ _01509_ VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10450_ _04354_ _04344_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09109_ _03019_ VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__buf_6
X_10381_ _04283_ Oset\[1\]\[9\] _03764_ _04286_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_75_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12120_ _05928_ _03874_ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12051_ _00639_ _00572_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11002_ _03685_ _04050_ _04903_ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__o21ai_1
X_12953_ clknet_3_5__leaf_clk _00396_ VGND VGND VPWR VPWR result_reg_set\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11904_ _02118_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12884_ clknet_leaf_23_clk _00327_ VGND VGND VPWR VPWR result_reg_Rshift\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_86_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
X_11835_ _05701_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__buf_4
X_11766_ _05628_ _04826_ _05653_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__o21ai_1
X_10717_ _03023_ Oset\[0\]\[10\] VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__nand2_1
X_11697_ H\[2\]\[15\] _04856_ _05596_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10648_ _02163_ _04552_ _02796_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_11_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10579_ _03770_ _04483_ _01156_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12318_ _06077_ _06078_ _02125_ VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12249_ _06033_ _00689_ VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06810_ _00930_ _00935_ _00608_ VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__mux2_1
X_07790_ _01447_ _01682_ VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06741_ net13 _00600_ _00739_ VGND VGND VPWR VPWR _00870_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09460_ _03366_ _03369_ VGND VGND VPWR VPWR _03370_ sky130_fd_sc_hd__nand2_1
X_06672_ _00785_ _00725_ _00802_ VGND VGND VPWR VPWR _00803_ sky130_fd_sc_hd__o21a_1
X_08411_ _02311_ _02318_ _02140_ _02326_ _02334_ VGND VGND VPWR VPWR _02335_ sky130_fd_sc_hd__o221ai_4
Xclkbuf_leaf_16_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09391_ _02947_ _02237_ _02904_ VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08342_ _02241_ Qset\[3\]\[5\] VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__nand2_1
X_08273_ Oset\[3\]\[2\] _02129_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__nor2_1
X_07224_ result_reg_set\[3\] VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07155_ _01238_ _00670_ VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__nand2_1
X_07086_ _00570_ Him _00573_ VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__or3_2
XFILLER_0_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07988_ _02006_ VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__clkbuf_1
X_06939_ result_reg_mul\[14\] VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__inv_2
X_09727_ Qset\[3\]\[7\] _03341_ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09658_ _03110_ _00556_ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09589_ _02992_ VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__buf_6
X_08609_ _02523_ Qset\[2\]\[0\] VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__nand2_1
X_11620_ _05341_ _04974_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11551_ _05437_ _05451_ VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_25_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10502_ _04407_ _04196_ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11482_ _04854_ _04460_ VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__nand2_1
X_10433_ _04194_ _04157_ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10364_ _03049_ _02735_ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__nor2_2
X_12103_ _01578_ _03072_ _03647_ VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__or3_1
X_10295_ _03506_ _03614_ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__nand2_1
X_12034_ _05844_ _05807_ _05857_ _05860_ VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__o211a_1
X_12936_ clknet_leaf_22_clk _00379_ VGND VGND VPWR VPWR result_reg_not\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12867_ clknet_leaf_23_clk _00310_ VGND VGND VPWR VPWR result_reg_Lshift\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ result_reg_mul\[10\] _05669_ _05682_ VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12798_ clknet_leaf_40_clk _00241_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11749_ _05642_ VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_5_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
X_08960_ _02871_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08891_ _02787_ Oset\[2\]\[2\] VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__nand2_1
X_07911_ _01951_ VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__clkbuf_1
X_07842_ _01893_ result_reg_mac\[13\] _01540_ VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__mux2_1
X_07773_ _01586_ result_reg_sub\[10\] VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__nand2_1
X_09512_ H\[3\]\[5\] _03033_ _03026_ VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__a21o_1
X_06724_ _00848_ _00853_ VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__nand2_4
XFILLER_0_91_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06655_ result_reg_set\[4\] VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__inv_2
X_09443_ _03351_ _03318_ _03319_ VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__nand3b_1
X_09374_ _03282_ _03284_ VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__nand2_1
X_06586_ _00707_ _00619_ _00719_ VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08325_ _02248_ _02249_ _02250_ _02251_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_50_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08256_ H\[2\]\[1\] VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_22_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07207_ _00726_ _01289_ _01181_ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__mux2_1
X_08187_ _02118_ CMD_addition VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07138_ _01220_ _01222_ VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07069_ _01153_ VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__buf_4
X_10080_ _03986_ _03983_ VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_58_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10982_ _04729_ Oset\[3\]\[12\] _04045_ VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_83_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12721_ clknet_leaf_33_clk _00164_ VGND VGND VPWR VPWR Oset\[1\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_12652_ clknet_leaf_37_clk _00102_ VGND VGND VPWR VPWR H\[3\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11603_ _04076_ _05335_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12583_ clknet_leaf_40_clk _00033_ VGND VGND VPWR VPWR Qset\[0\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11534_ _05196_ _05190_ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__nand2_1
X_11465_ _05364_ _05235_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10416_ _04320_ _04321_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_94_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11396_ _05296_ _03746_ _05297_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__nand3_2
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10347_ _03812_ _03814_ _04253_ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10278_ _04184_ _04151_ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12017_ _05763_ _05848_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12919_ clknet_leaf_31_clk _00362_ VGND VGND VPWR VPWR result_reg_or\[6\] sky130_fd_sc_hd__dfxtp_1
X_06440_ _00569_ _00574_ VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06371_ _00508_ _00509_ _06285_ VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__o21ai_1
X_08110_ _02071_ VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09090_ _02611_ VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__buf_6
X_08041_ Oset\[1\]\[14\] _01508_ _02018_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09992_ _03898_ VGND VGND VPWR VPWR _03899_ sky130_fd_sc_hd__buf_4
X_08943_ _02854_ _02833_ _02834_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__nand3b_1
X_08874_ _02522_ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__buf_6
X_07825_ result_reg_not\[12\] _01633_ _01877_ VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__a21o_1
X_07756_ _00930_ _01560_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__or2_1
X_06707_ _00829_ _00566_ _00732_ _00699_ VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_55_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07687_ _01559_ VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09426_ _03333_ _03335_ _02551_ VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__nand3_1
X_06638_ result_reg_sub\[3\] VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06569_ result_reg_add\[1\] VGND VGND VPWR VPWR _00703_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09357_ _03265_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08308_ _02230_ _02234_ _02143_ _02235_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__a211o_1
X_09288_ _03195_ _03198_ VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08239_ _02169_ VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11250_ _02469_ _04832_ _04835_ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10201_ _00589_ _04107_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__or2_2
X_11181_ _05081_ _05062_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__nand2_1
X_10132_ _04030_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__inv_2
X_10063_ _03968_ _03969_ VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12704_ clknet_leaf_3_clk _00009_ VGND VGND VPWR VPWR current_state\[2\] sky130_fd_sc_hd__dfxtp_4
X_10965_ _04865_ _04866_ _04867_ _04862_ _00647_ VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__a221o_1
X_10896_ H\[1\]\[11\] _03793_ _03798_ _04799_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__a211o_1
XFILLER_0_72_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12635_ clknet_leaf_38_clk _00085_ VGND VGND VPWR VPWR Oset\[3\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12566_ clknet_leaf_38_clk _00016_ VGND VGND VPWR VPWR next_PC\[2\] sky130_fd_sc_hd__dfxtp_1
X_11517_ _05416_ _05210_ VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12497_ _06214_ _01532_ VGND VGND VPWR VPWR _06215_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11448_ _05346_ _05347_ _05348_ _04859_ _00621_ VGND VGND VPWR VPWR _05349_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11379_ _05278_ _05279_ VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07610_ _01608_ _00755_ VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__nand2_1
X_08590_ _02502_ _02505_ VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__nand2_2
X_07541_ _01601_ _01604_ _01605_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__and3_2
X_07472_ _01536_ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__clkbuf_4
X_06423_ _00557_ current_state\[5\] VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09211_ _02525_ _03117_ _03119_ _03121_ VGND VGND VPWR VPWR _03122_ sky130_fd_sc_hd__o31ai_4
XTAP_TAPCELL_ROW_60_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06354_ _00491_ next_PC\[4\] VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__nand2_1
X_09142_ _02874_ _02312_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_32_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09073_ _02983_ _02981_ _02982_ VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__nand3_1
XFILLER_0_4_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08024_ _02025_ VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09975_ _03878_ _03881_ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__nand2_1
X_08926_ H\[3\]\[2\] _02836_ _02837_ _02838_ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__a211o_1
XFILLER_0_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08857_ _02766_ _02769_ _02551_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__nand3_1
X_07808_ _01016_ _01007_ _01544_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08788_ Oreg3 _02696_ _00626_ _02701_ VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__o211a_1
X_07739_ _01594_ _01788_ _01795_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10750_ _04652_ _04650_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10681_ _04575_ _04585_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__xnor2_1
X_09409_ _03316_ _03310_ _03313_ VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__nand3_1
X_12420_ _06256_ _06105_ VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__nand2_1
X_12351_ net22 net21 VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12282_ _00577_ _02119_ _02120_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__and3_1
X_11302_ _04952_ _04947_ VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__nand2_1
X_11233_ _05132_ _02649_ _05133_ _05135_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_73_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11164_ _03506_ _03110_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__nand2_1
X_11095_ _04996_ _04997_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__and2b_1
X_10115_ _04020_ _04012_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__nand2_1
X_10046_ _03952_ _03904_ VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11997_ _05834_ _05771_ VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_82_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10948_ _02442_ _00585_ _03768_ VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10879_ _04781_ _04782_ _04778_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__nand3_1
XFILLER_0_42_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12618_ clknet_leaf_34_clk _00068_ VGND VGND VPWR VPWR Qset\[2\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12549_ _06245_ VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_91_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1 _00073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06972_ result_reg_set\[15\] VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__inv_2
X_09760_ _03666_ _03519_ _03607_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__nand3b_1
X_09691_ _03598_ _03599_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__or2_2
X_08711_ _00001_ VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__inv_2
X_08642_ _01959_ _01154_ _02556_ VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_1_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08573_ H\[3\]\[14\] VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_65_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07524_ _01588_ VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07455_ _01276_ _01511_ _01523_ _01524_ VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__a22o_1
X_06406_ _00540_ VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__clkbuf_4
X_07386_ result_reg_and\[12\] _01299_ VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06337_ _00480_ VGND VGND VPWR VPWR _00481_ sky130_fd_sc_hd__inv_2
X_09125_ _03022_ Qset\[2\]\[4\] VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__nand2_1
X_09056_ Qset\[3\]\[3\] _02836_ _02837_ VGND VGND VPWR VPWR _02968_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08007_ Oset\[0\]\[14\] _01508_ _02000_ VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09958_ _02420_ _02544_ VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__nand2_1
X_08909_ _02687_ _02821_ VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__nand2_1
X_09889_ _03793_ _02346_ VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__nor2_1
X_11920_ _00591_ _05767_ VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__nor2_1
X_11851_ _05714_ VGND VGND VPWR VPWR _00295_ sky130_fd_sc_hd__inv_2
X_11782_ _05665_ VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__inv_2
X_10802_ _04705_ _04648_ VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__nand2_1
X_10733_ _04637_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10664_ _04567_ _04568_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__nand2_1
X_12403_ _06135_ _06253_ _06267_ _06143_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__a211o_1
X_10595_ _04463_ _04467_ _04464_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__nand3_1
X_12334_ _06087_ VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__clkbuf_1
X_12265_ _06039_ _05813_ _06013_ _06043_ VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12196_ _05960_ _05991_ VGND VGND VPWR VPWR _05992_ sky130_fd_sc_hd__nand2_1
X_11216_ _04830_ _04896_ _03283_ _05116_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__o211ai_1
Xoutput60 net60 VGND VGND VPWR VPWR data_out[6] sky130_fd_sc_hd__buf_1
X_11147_ _05048_ _05049_ VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__nand2_1
Xoutput71 net71 VGND VGND VPWR VPWR instruction_address[6] sky130_fd_sc_hd__buf_1
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11078_ _04980_ _03079_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__nand2_1
X_10029_ _03933_ _03934_ VGND VGND VPWR VPWR _03936_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07240_ net11 _01193_ VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__nor2_1
X_07171_ _01193_ VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_14_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09812_ Qset\[1\]\[7\] _03033_ VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06955_ result_reg_Lshift\[14\] VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__inv_2
X_09743_ _03650_ _02334_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__nand2_4
X_06886_ result_reg_sub\[12\] _00541_ _01008_ VGND VGND VPWR VPWR _01009_ sky130_fd_sc_hd__o21ai_1
X_09674_ _03021_ Qset\[0\]\[6\] VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08625_ _02539_ VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__buf_4
X_08556_ _02311_ _02458_ _02139_ _02466_ _02473_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_76_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07507_ _01196_ _01571_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__nand2_4
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08487_ _02328_ _02406_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__nor2_1
X_07438_ Oset\[3\]\[14\] _01508_ _01249_ VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07369_ _00991_ _01267_ _01263_ _01442_ VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09108_ _03018_ _02264_ VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__nand2_2
XFILLER_0_60_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10380_ _04283_ _02368_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_75_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09039_ _02916_ _02950_ VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__nand2_1
X_12050_ _05844_ _05841_ _05857_ _05869_ VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__o211a_1
X_11001_ _03685_ _04050_ _04903_ VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__or3_1
XFILLER_0_99_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12952_ clknet_leaf_15_clk _00395_ VGND VGND VPWR VPWR result_reg_set\[7\] sky130_fd_sc_hd__dfxtp_1
X_11903_ _01158_ _02807_ _02817_ _05749_ _05752_ VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__a221o_2
X_12883_ clknet_leaf_23_clk _00326_ VGND VGND VPWR VPWR result_reg_Rshift\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_86_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _05667_ _04830_ _00528_ VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11765_ _05628_ _00991_ _02650_ VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11696_ H\[3\]\[15\] _04858_ _04859_ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__a21o_1
X_10716_ _04617_ _04618_ _03794_ _04619_ _04620_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__a32o_1
X_10647_ _04549_ _04551_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__nand2_2
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10578_ _04479_ _04480_ _04481_ _04482_ VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__o22a_2
XTAP_TAPCELL_ROW_97_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12317_ _05766_ _06059_ VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12248_ _06032_ _05748_ _06013_ _06034_ VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__o211a_1
X_12179_ _05903_ _05902_ VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06740_ result_reg_set\[6\] _00615_ _00696_ _00868_ VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06671_ _00794_ _00619_ _00629_ _00801_ VGND VGND VPWR VPWR _00802_ sky130_fd_sc_hd__a211o_1
XFILLER_0_64_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08410_ _02331_ _02333_ _01552_ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__a21o_2
X_09390_ _02954_ _03268_ _03264_ VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_58_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08341_ _02230_ Qset\[2\]\[5\] VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08272_ _02197_ _02200_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07223_ result_reg_or\[3\] _01199_ VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07154_ R2\[1\] _01238_ VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07085_ result_reg_set\[0\] VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07987_ Oset\[0\]\[4\] _01332_ _02001_ VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__mux2_1
X_06938_ result_reg_sub\[14\] _00541_ _01058_ VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__o21ai_2
X_09726_ _02318_ _02162_ VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__nand2_1
X_06869_ _00985_ _00992_ _00732_ VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__mux2_1
X_09657_ _03536_ _00623_ _03565_ VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__nand3_1
XFILLER_0_96_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09588_ _03341_ H\[2\]\[6\] VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__nand2_1
X_08608_ _02522_ VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__buf_4
X_08539_ _02397_ Qset\[1\]\[13\] _02378_ _02456_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__a211o_1
XFILLER_0_64_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11550_ _05449_ _05450_ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10501_ _04401_ _04402_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11481_ _04458_ _05157_ VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10432_ _04337_ _03746_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10363_ _04268_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12102_ _01359_ _05873_ _05913_ _05914_ _02650_ VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__a221oi_1
X_12033_ _05844_ _00922_ VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__nand2_1
X_10294_ _04200_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__inv_2
X_12935_ clknet_leaf_22_clk _00378_ VGND VGND VPWR VPWR result_reg_not\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12866_ clknet_leaf_24_clk _00309_ VGND VGND VPWR VPWR result_reg_Lshift\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_44_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ _05690_ VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__inv_2
X_12797_ clknet_leaf_40_clk _00240_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_99_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _00841_ _05631_ _05634_ _05641_ VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__a211o_1
XFILLER_0_83_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11679_ _02897_ _05158_ VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08890_ _02802_ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__inv_2
X_07910_ Oset\[2\]\[8\] _01403_ _01942_ VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__mux2_1
X_07841_ _01593_ _01886_ _01892_ VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07772_ _01581_ result_reg_add\[10\] VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__nand2_1
X_06723_ _00849_ _00655_ _00657_ _00852_ _00666_ VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__a221o_2
XFILLER_0_78_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09511_ _03349_ VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__buf_6
XFILLER_0_78_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06654_ result_reg_mac\[4\] VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__inv_2
X_09442_ _03320_ _03351_ VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__nand2_1
X_06585_ _00708_ _00709_ _00714_ _00718_ _00603_ VGND VGND VPWR VPWR _00719_ sky130_fd_sc_hd__o221a_1
XFILLER_0_59_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09373_ _03277_ _03278_ _03283_ VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__nand3_1
XFILLER_0_19_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08324_ _02248_ Oset\[3\]\[4\] VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08255_ _02181_ _02184_ VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__nand2_1
X_07206_ _00727_ _01288_ _01176_ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__mux2_1
X_08186_ shift.left VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__buf_4
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07137_ _00681_ _01190_ _01221_ VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07068_ _00583_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10981_ _04881_ _02436_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__nor2_1
X_09709_ _03616_ _03421_ _03462_ VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__nand3_1
X_12720_ clknet_leaf_38_clk _00163_ VGND VGND VPWR VPWR Oset\[1\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_83_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12651_ clknet_leaf_32_clk _00101_ VGND VGND VPWR VPWR H\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11602_ _04302_ _02503_ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12582_ clknet_leaf_40_clk _00032_ VGND VGND VPWR VPWR Qset\[0\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11533_ _05205_ _05201_ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11464_ _05235_ _05364_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10415_ _03411_ VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11395_ _05114_ _05294_ _05230_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10346_ _04251_ _04252_ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__nand2_1
X_10277_ _04142_ _04143_ _04150_ VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__a21o_1
X_12016_ result_reg_Rshift\[1\] _05848_ _05808_ _05849_ VGND VGND VPWR VPWR _00325_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12918_ clknet_leaf_16_clk _00361_ VGND VGND VPWR VPWR result_reg_or\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ clknet_leaf_10_clk _00292_ VGND VGND VPWR VPWR result_reg_mac\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06370_ _00501_ _00506_ VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__and2_1
X_08040_ _02033_ VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09991_ _03835_ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08942_ _02835_ _02854_ VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08873_ _02785_ _02577_ VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__and2_1
X_07824_ result_reg_Rshift\[12\] _01672_ _01601_ _01876_ VGND VGND VPWR VPWR _01877_
+ sky130_fd_sc_hd__o211a_1
X_07755_ _01809_ _01653_ _01810_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__a21o_1
X_07686_ _01353_ _01682_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__or2_1
X_06706_ _00818_ _00819_ _00835_ VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_55_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06637_ _00553_ result_reg_or\[3\] VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__or2b_1
XFILLER_0_94_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09425_ _02992_ _02277_ _03004_ _03334_ VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__o211ai_2
X_06568_ result_reg_sub\[1\] VGND VGND VPWR VPWR _00702_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09356_ _03266_ _02954_ VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__nand2_1
X_06499_ _00529_ VGND VGND VPWR VPWR _00634_ sky130_fd_sc_hd__buf_2
X_08307_ H\[1\]\[3\] _02230_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__nor2_1
X_09287_ _03196_ _03197_ VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08238_ _02168_ VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__clkbuf_4
X_08169_ R2\[1\] _02100_ _02105_ _02108_ VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__o211a_1
X_10200_ _04042_ _04103_ _04104_ _04106_ VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_42_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11180_ _05082_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__inv_2
X_10131_ _04034_ _04035_ _04037_ VGND VGND VPWR VPWR _04038_ sky130_fd_sc_hd__nand3_1
X_10062_ _03967_ _03962_ VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12703_ clknet_leaf_3_clk _00008_ VGND VGND VPWR VPWR current_state\[1\] sky130_fd_sc_hd__dfxtp_1
X_10964_ _02436_ _04838_ _04858_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10895_ _03793_ _03861_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__nor2_1
X_12634_ clknet_leaf_37_clk _00084_ VGND VGND VPWR VPWR Oset\[3\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12565_ clknet_leaf_39_clk _00015_ VGND VGND VPWR VPWR next_PC\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11516_ _05210_ _05416_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12496_ R3\[0\] net17 current_state\[2\] VGND VGND VPWR VPWR _06214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11447_ _02479_ _04053_ _03793_ VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11378_ _05254_ _05278_ _05279_ VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__nand3b_1
X_10329_ _03229_ _03232_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07540_ _01555_ _00640_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07471_ Hreg3 VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__buf_4
X_06422_ CMD_multiplication VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09210_ _02562_ Oset\[3\]\[5\] _02800_ _03120_ VGND VGND VPWR VPWR _03121_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_101_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06353_ _00489_ _00475_ _00494_ next_PC\[3\] _00478_ VGND VGND VPWR VPWR _00017_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09141_ _03051_ _02738_ VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_60_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09072_ _02981_ _02982_ _02983_ VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08023_ Oset\[1\]\[5\] _01349_ _02019_ VGND VGND VPWR VPWR _02025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09974_ _03879_ _03880_ VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__nand2_1
X_08925_ _02688_ _02207_ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08856_ _02767_ _02590_ _02768_ VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__nand3_2
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07807_ _01860_ VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__clkbuf_1
X_08787_ _02698_ _02700_ _00646_ VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__a21o_1
X_07738_ _01792_ _01572_ _01793_ _01568_ _01794_ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__a311o_1
XFILLER_0_67_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07669_ _01579_ result_reg_sub\[5\] VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_80_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10680_ _04583_ _04584_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__and2b_1
X_09408_ _03314_ _03317_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__nand2_1
X_09339_ _03244_ _03249_ VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12350_ net24 net25 VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__nor2_1
X_12281_ _02099_ _02165_ VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__and2_1
X_11301_ _05202_ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11232_ result_reg_add\[12\] _02649_ _05134_ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_91_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11163_ _03690_ _05065_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__or2_1
X_10114_ _04012_ _04020_ VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__or2_1
X_11094_ _04995_ _04983_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__nand2_1
X_10045_ _03917_ _03913_ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11996_ _05821_ _05833_ _05754_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10947_ _03781_ _04842_ _00584_ _04849_ VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10878_ _04571_ _04568_ _04758_ VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__nand3_1
X_12617_ clknet_leaf_35_clk _00067_ VGND VGND VPWR VPWR Qset\[2\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12548_ _00979_ Qset\[3\]\[10\] _06233_ VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12479_ _06267_ _00582_ _06202_ _06204_ _05775_ VGND VGND VPWR VPWR _06205_ sky130_fd_sc_hd__a221o_1
XANTENNA_2 _00473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06971_ _01089_ _01090_ _00835_ VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__a21o_1
X_09690_ _03597_ _03444_ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__and2_1
X_08710_ _02624_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__clkbuf_4
X_08641_ _02555_ VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_1_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08572_ _02485_ _02488_ VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_65_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07523_ _00559_ _01571_ VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__nand2_1
X_07454_ _01082_ _01275_ _01160_ VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06405_ _00539_ VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__buf_2
XFILLER_0_91_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07385_ result_reg_not\[12\] _01457_ _01167_ VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06336_ next_PC\[1\] next_PC\[0\] VGND VGND VPWR VPWR _00480_ sky130_fd_sc_hd__nand2_1
X_09124_ Qset\[3\]\[4\] _03025_ _03027_ VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09055_ H\[1\]\[3\] _02836_ _02840_ _02966_ VGND VGND VPWR VPWR _02967_ sky130_fd_sc_hd__a211o_1
X_08006_ _02015_ VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_77_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09957_ _02561_ H\[2\]\[11\] _02727_ VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__o21a_1
X_08908_ _02819_ _02820_ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__nand2_4
XFILLER_0_99_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09888_ _03794_ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__clkbuf_4
X_08839_ _02752_ VGND VGND VPWR VPWR _00245_ sky130_fd_sc_hd__inv_2
X_11850_ _00761_ _05707_ _05710_ _05713_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__a211o_1
XFILLER_0_86_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11781_ _05663_ _05664_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10801_ _04701_ _04703_ _04704_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__nand3_1
XFILLER_0_67_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10732_ _04635_ _04636_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10663_ _04564_ _04566_ _04565_ VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__nand3_2
X_12402_ _06139_ _06142_ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10594_ _04496_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12333_ _01529_ _01532_ VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__and2_1
X_12264_ result_reg_not\[8\] _06031_ VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__or2b_1
X_11215_ _05117_ _03281_ VGND VGND VPWR VPWR _05118_ sky130_fd_sc_hd__nand2_1
X_12195_ _05789_ _03639_ _05907_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__a21o_1
Xoutput61 net61 VGND VGND VPWR VPWR data_out[7] sky130_fd_sc_hd__buf_1
Xoutput50 net50 VGND VGND VPWR VPWR data_out[11] sky130_fd_sc_hd__buf_1
X_11146_ _05046_ _05044_ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__or2b_1
Xoutput72 net72 VGND VGND VPWR VPWR instruction_address[7] sky130_fd_sc_hd__buf_1
X_11077_ _04095_ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__inv_2
X_10028_ _03926_ _03933_ _03934_ VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_62_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11979_ result_reg_Lshift\[10\] _05743_ _05808_ _05819_ VGND VGND VPWR VPWR _00318_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07170_ _01190_ VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_8 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09811_ _03021_ Qset\[0\]\[7\] VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__nand2_1
X_09742_ _03649_ _01552_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__nand2_1
X_06954_ result_reg_not\[14\] VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06885_ _00540_ _01007_ _00534_ VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__a21oi_1
X_09673_ _03578_ _03579_ _03026_ _03580_ _03581_ VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__a32o_1
X_08624_ Oreg3 Oreg2 VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__nor2_4
X_08555_ _02468_ _02472_ _01554_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__a21o_1
X_07506_ Hreg2 VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__buf_4
XFILLER_0_76_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08486_ Qset\[2\]\[11\] VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07437_ _01161_ _01493_ _01507_ VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_76_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07368_ result_reg_add\[11\] _01267_ VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06319_ LC\[6\] _06279_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09107_ _03017_ _01552_ VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__nand2_2
X_07299_ result_reg_and\[7\] _01207_ _01261_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09038_ _02578_ _02949_ VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__nor2_1
X_11000_ _04766_ _04901_ _04902_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__o21ai_1
X_12951_ clknet_leaf_15_clk _00394_ VGND VGND VPWR VPWR result_reg_set\[6\] sky130_fd_sc_hd__dfxtp_1
X_12882_ clknet_leaf_24_clk _00325_ VGND VGND VPWR VPWR result_reg_Rshift\[1\] sky130_fd_sc_hd__dfxtp_1
X_11902_ _00591_ _05751_ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ result_reg_mul\[15\] _05670_ _05672_ _05700_ VGND VGND VPWR VPWR _00291_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11764_ _05652_ VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11695_ _05593_ _05594_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10715_ _03023_ Qset\[2\]\[10\] VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10646_ _04105_ Qset\[1\]\[10\] _04042_ _04550_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__a211o_1
XFILLER_0_36_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10577_ Oset\[1\]\[10\] _03773_ _03761_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_97_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12316_ _00956_ _06058_ VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12247_ _06033_ _00652_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__nand2_1
X_12178_ result_reg_or\[3\] _05959_ _05976_ _05977_ _05940_ VGND VGND VPWR VPWR _00359_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11129_ _04978_ _05031_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__nand2_1
X_06670_ _00795_ _00709_ _00739_ _00800_ VGND VGND VPWR VPWR _00801_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08340_ _02266_ VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__clkbuf_1
X_08271_ _02198_ _02135_ _02199_ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__nand3_1
X_07222_ _01300_ _01303_ _01271_ VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07153_ _00634_ _01231_ _01235_ _01236_ _01237_ VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_42_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07084_ result_reg_not\[0\] _01166_ _01168_ VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07986_ _02005_ VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__clkbuf_1
X_06937_ _00740_ _01057_ _00535_ VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__a21oi_1
X_09725_ _02540_ _03632_ _01155_ VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__o21ai_1
X_09656_ _03564_ _03233_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__nand2_1
X_06868_ _00991_ _00982_ _00730_ VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__mux2_1
X_08607_ _00006_ VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__clkinv_4
X_06799_ result_reg_not\[8\] _00921_ _00925_ _00664_ VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09587_ _03495_ _02556_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08538_ _02397_ _02455_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08469_ _02386_ _02389_ VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__nand2_2
XFILLER_0_37_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10500_ _04404_ _00831_ _04405_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__nand3_1
X_11480_ _05093_ _05260_ _05265_ VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10431_ _04335_ _04336_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10362_ _04267_ _04202_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12101_ _05892_ _03489_ _05783_ _05878_ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__o31a_1
XFILLER_0_20_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10293_ _03624_ _03621_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__nand2_1
X_12032_ _05844_ _05801_ _05857_ _05859_ VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12934_ clknet_leaf_22_clk _00377_ VGND VGND VPWR VPWR result_reg_not\[5\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12865_ clknet_leaf_20_clk _00308_ VGND VGND VPWR VPWR result_reg_Lshift\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11816_ _04408_ _04409_ _05677_ _05689_ VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__a31o_1
X_12796_ clknet_leaf_41_clk _00239_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11747_ _05627_ _03449_ VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11678_ _04854_ _02895_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10629_ _04533_ _04362_ _04360_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07840_ _01041_ _01574_ _01890_ _01891_ _01569_ VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__a221o_1
X_07771_ _01823_ _01658_ _01824_ _01825_ VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06722_ result_reg_Rshift\[5\] _00753_ _00851_ VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__o21ai_1
X_09510_ _03418_ _00536_ _03419_ VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09441_ _03350_ _03258_ VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__nor2_1
X_06653_ _00784_ VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__clkbuf_1
X_06584_ _00715_ _00717_ _00560_ VGND VGND VPWR VPWR _00718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09372_ _03281_ VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08323_ _02143_ VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08254_ _02127_ _02182_ _02135_ _02183_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__o211ai_1
X_07205_ _00728_ _00729_ _01173_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__mux2_1
X_08185_ _02116_ _02117_ VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__nor2_1
X_07136_ _01190_ R0\[0\] VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07067_ _01152_ VGND VGND VPWR VPWR _00073_ sky130_fd_sc_hd__buf_1
XFILLER_0_30_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07969_ LC\[7\] _01992_ _01993_ _01994_ VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__a22o_1
X_09708_ _03020_ _03614_ VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_58_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10980_ _03152_ Oset\[0\]\[12\] _04042_ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__a21oi_1
X_09639_ _03387_ _03545_ _03547_ VGND VGND VPWR VPWR _03548_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12650_ clknet_leaf_41_clk _00100_ VGND VGND VPWR VPWR H\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11601_ _02506_ _02163_ _03781_ VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12581_ clknet_leaf_43_clk _00031_ VGND VGND VPWR VPWR Qset\[0\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11532_ _05431_ _05432_ _03751_ VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__nand3_1
X_11463_ _05063_ _03110_ VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_21_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10414_ _04318_ _04319_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11394_ _05231_ _05295_ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_94_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10345_ _00710_ _03835_ _00831_ _04249_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__o211ai_1
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10276_ _04010_ _04182_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__nand2_1
X_12015_ _05756_ _05848_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12917_ clknet_leaf_17_clk _00360_ VGND VGND VPWR VPWR result_reg_or\[4\] sky130_fd_sc_hd__dfxtp_1
X_12848_ clknet_leaf_7_clk _00291_ VGND VGND VPWR VPWR result_reg_mul\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ clknet_leaf_24_clk _00222_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09990_ _03049_ VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__clkbuf_4
X_08941_ _00622_ _02785_ _02853_ VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08872_ _02784_ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__buf_6
X_07823_ _01716_ _01025_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__nand2_1
X_07754_ result_reg_mul\[9\] _01548_ _01656_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07685_ _01742_ _01549_ _01743_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__a21o_1
X_06705_ _00635_ _00824_ _00828_ _00830_ _00834_ VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__o2111ai_4
XTAP_TAPCELL_ROW_55_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06636_ _00764_ _00562_ _00766_ _00767_ VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__a31o_1
X_09424_ _03001_ Oset\[1\]\[5\] VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06567_ result_reg_mul\[1\] VGND VGND VPWR VPWR _00701_ sky130_fd_sc_hd__inv_2
X_09355_ _03264_ _03265_ VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__nand2b_1
X_06498_ _00631_ _00632_ VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__nor2_2
X_08306_ H\[0\]\[3\] VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__inv_2
X_09286_ _03194_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__inv_2
X_08237_ _00635_ _02166_ _02167_ VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__or3_2
XFILLER_0_34_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_08168_ _02102_ _02103_ net41 VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__a21o_1
X_07119_ _01200_ _00533_ VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__nor2_4
X_08099_ _01801_ H\[1\]\[8\] _02057_ VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10130_ _03983_ _04036_ _04007_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10061_ _03962_ _03967_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__or2_1
X_10963_ _04856_ Oset\[0\]\[12\] _04862_ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__a21oi_1
X_12702_ clknet_leaf_3_clk net35 VGND VGND VPWR VPWR current_state\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10894_ H\[2\]\[11\] _04415_ _04797_ VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__a21o_1
X_12633_ clknet_leaf_40_clk _00083_ VGND VGND VPWR VPWR Oset\[3\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_12564_ clknet_leaf_39_clk _00014_ VGND VGND VPWR VPWR next_PC\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11515_ _04854_ _04955_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12495_ _06213_ VGND VGND VPWR VPWR _00440_ sky130_fd_sc_hd__clkbuf_1
X_11446_ Qset\[3\]\[14\] _04857_ _04859_ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11377_ _05277_ _05274_ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10328_ _04233_ _04234_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10259_ _04165_ _03944_ VGND VGND VPWR VPWR _04166_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07470_ _01535_ VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__clkbuf_1
X_06421_ _00549_ VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__buf_4
XFILLER_0_29_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06352_ _06285_ _00493_ VGND VGND VPWR VPWR _00494_ sky130_fd_sc_hd__nand2_1
X_09140_ _03048_ _03050_ VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_60_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09071_ _02859_ _02856_ VGND VGND VPWR VPWR _02983_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08022_ _02024_ VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09973_ _02687_ _03868_ VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__nand2_1
X_08924_ _02626_ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__clkbuf_4
X_08855_ _02579_ Oset\[1\]\[2\] VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_68_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08786_ Oset\[1\]\[1\] _02625_ _00001_ _02699_ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__a211o_1
X_07806_ _01859_ H\[3\]\[11\] _01628_ VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__mux2_1
X_07737_ result_reg_or\[8\] _01595_ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07668_ _01580_ result_reg_add\[5\] VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_80_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06619_ result_reg_not\[2\] VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__inv_2
X_07599_ _01586_ result_reg_sub\[2\] VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__nand2_1
X_09407_ _03316_ VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__inv_2
X_09338_ _03246_ _03247_ _03248_ VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__nand3_1
XFILLER_0_35_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11300_ _05200_ _05201_ VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09269_ _03179_ _03107_ VGND VGND VPWR VPWR _03180_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12280_ _06031_ _05838_ _06044_ _06051_ VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__o211a_1
X_11231_ _00472_ VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11162_ _03505_ _03076_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10113_ _04018_ _04019_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__nand2_1
X_11093_ _04983_ _04995_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__nor2_1
X_10044_ _03948_ _03950_ VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11995_ _04071_ _05749_ _04064_ _05745_ _05832_ VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__a221o_2
XFILLER_0_58_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10946_ _02162_ _02435_ _03781_ _04848_ VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_85_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10877_ _04724_ _04757_ VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_100_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12616_ clknet_leaf_35_clk _00066_ VGND VGND VPWR VPWR Qset\[2\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12547_ _06244_ VGND VGND VPWR VPWR _00461_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12478_ _06130_ _06186_ _06139_ _06171_ _06203_ VGND VGND VPWR VPWR _06204_ sky130_fd_sc_hd__o221a_1
XFILLER_0_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_3 _00498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11429_ _02482_ _02163_ _03781_ VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__a21o_1
X_06970_ _00714_ result_reg_or\[15\] VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__nand2_1
X_08640_ Hreg3 Hreg2 VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_1_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08571_ _02470_ Oset\[1\]\[14\] _02444_ _02487_ VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_65_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_46_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07522_ _01586_ result_reg_sub\[0\] VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__nand2_1
X_07453_ _01192_ _01516_ _01517_ _01220_ _01522_ VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__a311o_1
XFILLER_0_76_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06404_ _00538_ _00526_ VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07384_ result_reg_Lshift\[12\] result_reg_Rshift\[12\] _01164_ VGND VGND VPWR VPWR
+ _01457_ sky130_fd_sc_hd__mux2_1
X_09123_ Qset\[1\]\[4\] _03033_ VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__nand2_1
X_06335_ R3\[1\] _06285_ VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09054_ _02836_ _02234_ VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08005_ Oset\[0\]\[13\] _01490_ _02000_ VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09956_ _02423_ _02528_ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__nand2_1
X_08907_ R2\[0\] _00587_ VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__nand2_1
X_09887_ _03027_ VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__clkbuf_4
X_08838_ _00703_ _02654_ _02650_ _02751_ VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__a211o_1
XFILLER_0_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_37_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
X_08769_ _02682_ _02571_ VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__nand2_1
X_11780_ _05628_ _01093_ _02650_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10800_ _04455_ _04506_ _04697_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__nand3_1
XFILLER_0_79_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10731_ _04434_ _04631_ _04633_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__nand3b_1
X_12401_ _06141_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__inv_2
X_10662_ _04564_ _04565_ _04566_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__a21o_1
X_10593_ _04465_ _04469_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12332_ _06086_ VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__clkbuf_1
X_12263_ _06039_ _05793_ _06013_ _06042_ VGND VGND VPWR VPWR _00379_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11214_ _04830_ _04896_ _05116_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput40 net40 VGND VGND VPWR VPWR data_address[2] sky130_fd_sc_hd__buf_1
X_12194_ result_reg_or\[6\] _05959_ _05988_ _05990_ _05940_ VGND VGND VPWR VPWR _00362_
+ sky130_fd_sc_hd__o221a_1
Xoutput51 net51 VGND VGND VPWR VPWR data_out[12] sky130_fd_sc_hd__buf_1
X_11145_ _05043_ _05047_ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__nand2_1
Xoutput73 net73 VGND VGND VPWR VPWR instruction_address[8] sky130_fd_sc_hd__clkbuf_1
Xoutput62 net62 VGND VGND VPWR VPWR data_out[8] sky130_fd_sc_hd__buf_1
X_11076_ _04959_ _04978_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__and2b_1
X_10027_ _03932_ _03927_ VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_28_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
X_11978_ _05818_ _05771_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_62_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10929_ _04283_ VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__buf_6
XFILLER_0_46_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09810_ _03714_ _03715_ _03027_ _03716_ _03717_ VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__a32o_1
X_06953_ _01056_ _00695_ _01065_ _01073_ _00644_ VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__a221o_1
X_09741_ _03643_ _03648_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__nand2_1
X_06884_ result_reg_add\[12\] VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__inv_2
X_09672_ _03021_ Oset\[2\]\[6\] VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_6_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_19_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_27_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08623_ _02531_ _02537_ VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__nand2_1
X_08554_ _02469_ _02470_ _02444_ _02471_ VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07505_ _01540_ VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08485_ _02405_ VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__clkbuf_1
X_07436_ _01498_ _01214_ _01505_ _01159_ _01506_ VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__a311o_1
XFILLER_0_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07367_ result_reg_and\[11\] _01299_ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06318_ _06278_ VGND VGND VPWR VPWR _06279_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09106_ _03010_ _03016_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07298_ _01375_ _01255_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__nand2_1
X_09037_ _02948_ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09939_ _03843_ _03845_ VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__nand2_2
X_12950_ clknet_leaf_1_clk _00393_ VGND VGND VPWR VPWR result_reg_set\[5\] sky130_fd_sc_hd__dfxtp_1
X_12881_ clknet_leaf_21_clk _00324_ VGND VGND VPWR VPWR result_reg_Rshift\[0\] sky130_fd_sc_hd__dfxtp_1
X_11901_ _05750_ VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _05554_ _05592_ _05673_ VGND VGND VPWR VPWR _05700_ sky130_fd_sc_hd__a21o_1
X_11763_ _00958_ _05631_ _05634_ _05651_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__a211o_1
XFILLER_0_67_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11694_ _04980_ _02096_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10714_ Qset\[3\]\[10\] _03791_ _03794_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10645_ _04105_ _02391_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_11_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12315_ _06075_ _06055_ _06066_ _06076_ VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__o211a_1
X_10576_ _04282_ Oset\[0\]\[10\] VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_97_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12246_ _06031_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__buf_2
X_12177_ _05904_ _02944_ _05898_ _05957_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__a211o_1
X_11128_ _04309_ _04975_ _04977_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_79_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11059_ _04881_ Qset\[1\]\[13\] _04042_ _04961_ VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_88_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08270_ _02127_ Qset\[1\]\[2\] VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07221_ _00765_ _01266_ _01299_ _01302_ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07152_ _00831_ _00833_ _06264_ _00634_ _01171_ VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__a2111o_1
X_07083_ _01167_ VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_8_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_74_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07985_ Oset\[0\]\[3\] _01314_ _02001_ VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__mux2_1
X_06936_ result_reg_add\[14\] VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__inv_2
X_09724_ _03629_ _03631_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__nand2_2
X_06867_ result_reg_sub\[11\] VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__inv_2
X_09655_ _03562_ _03563_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08606_ _02521_ VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06798_ _00924_ _00656_ VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09586_ _03493_ _03494_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08537_ Qset\[0\]\[13\] VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08468_ _02364_ Oset\[1\]\[10\] _02378_ _02388_ VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__a211o_1
XFILLER_0_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07419_ Oset\[3\]\[13\] _01490_ _01249_ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08399_ Oset\[0\]\[7\] VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__inv_2
X_10430_ _04333_ _04246_ _04334_ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__nand3_1
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10361_ _03651_ _03462_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__nand2_1
X_12100_ _01578_ _03102_ _03502_ _05912_ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__o31a_1
X_10292_ _03655_ _03625_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__and2_1
X_12031_ _05844_ _00900_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12933_ clknet_leaf_19_clk _00376_ VGND VGND VPWR VPWR result_reg_not\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12864_ clknet_leaf_10_clk _00307_ VGND VGND VPWR VPWR result_reg_mac\[15\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_44_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11815_ result_reg_mul\[9\] _05669_ _05682_ VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__o21ai_1
X_12795_ clknet_leaf_44_clk _00238_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11746_ _05640_ VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11677_ _05575_ _05576_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_24_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10628_ _04011_ _04027_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10559_ _04462_ _04459_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12229_ _05958_ _06018_ VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07770_ net2 _01746_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__nor2_1
X_06721_ _00754_ _00850_ VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09440_ _03349_ VGND VGND VPWR VPWR _03350_ sky130_fd_sc_hd__inv_2
X_06652_ _00783_ Qset\[0\]\[3\] _00687_ VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_96_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06583_ _00716_ _00701_ _00534_ VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__mux2_1
X_09371_ _03279_ _03281_ VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08322_ Oset\[2\]\[4\] VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__inv_2
X_08253_ _02127_ Oset\[1\]\[1\] VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__nand2_1
X_07204_ _00738_ _01208_ _01190_ _01286_ VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08184_ _02102_ _02103_ net36 VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07135_ _01214_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__inv_2
X_07066_ _01151_ _01149_ VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07968_ _01990_ _01960_ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__nand2_1
X_06919_ result_reg_or\[13\] VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__inv_2
X_09707_ _03612_ _03020_ _03614_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07899_ _01945_ VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__clkbuf_1
X_09638_ _03385_ _03546_ VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_83_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09569_ _02611_ _02299_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__nor2_1
X_11600_ _05499_ VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__inv_2
X_12580_ clknet_leaf_44_clk _00030_ VGND VGND VPWR VPWR Qset\[0\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11531_ _05430_ _05225_ _05222_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_92_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11462_ _04308_ _03745_ _03145_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_21_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11393_ _05294_ VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__inv_2
X_10413_ _04234_ _04261_ _04316_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10344_ _04250_ _02160_ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_94_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10275_ _03986_ _03983_ _04008_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__nand3_1
X_12014_ _05847_ VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__buf_2
X_12916_ clknet_leaf_15_clk _00359_ VGND VGND VPWR VPWR result_reg_or\[3\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_29_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ clknet_leaf_5_clk _00290_ VGND VGND VPWR VPWR result_reg_mul\[14\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_56_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12778_ clknet_leaf_25_clk _00221_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dfxtp_1
X_11729_ _05627_ VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__buf_6
XFILLER_0_56_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08940_ _01536_ _02839_ _02842_ _00548_ _02852_ VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__a311o_1
XFILLER_0_20_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08871_ _02783_ _02213_ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__nand2_2
X_07822_ _01874_ result_reg_mac\[12\] _01540_ VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07753_ _00932_ _00933_ _01544_ VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__mux2_1
X_07684_ result_reg_mul\[6\] _01679_ _01656_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__o21ai_1
X_06704_ _00832_ _00833_ _06264_ _00635_ _00829_ VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_55_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06635_ result_reg_and\[3\] _00743_ _00553_ VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__o21ai_1
X_09423_ _03001_ _02274_ _02991_ _03332_ VGND VGND VPWR VPWR _03333_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_35_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09354_ _03263_ _03237_ VGND VGND VPWR VPWR _03265_ sky130_fd_sc_hd__nand2_1
X_06566_ result_reg_set\[1\] VGND VGND VPWR VPWR _00700_ sky130_fd_sc_hd__inv_2
X_08305_ _02230_ _02231_ _02147_ _02232_ VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__a211o_1
XFILLER_0_74_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06497_ CMD_or CMD_multiplication _00578_ VGND VGND VPWR VPWR _00632_ sky130_fd_sc_hd__or3_4
X_09285_ _03191_ _03193_ VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__nor2_1
X_08236_ _02099_ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08167_ R2\[0\] _02100_ _02105_ _02107_ VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__o211a_1
X_07118_ result_reg_add\[0\] result_reg_sub\[0\] _01202_ VGND VGND VPWR VPWR _01203_
+ sky130_fd_sc_hd__mux2_1
X_08098_ _02065_ VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07049_ _01004_ Qset\[2\]\[11\] _01128_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10060_ _03964_ _03966_ VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10962_ Oset\[1\]\[12\] _04858_ VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__nand2_1
X_12701_ clknet_leaf_30_clk _00151_ VGND VGND VPWR VPWR Oset\[0\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_10893_ H\[3\]\[11\] _03793_ _03795_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__a21o_1
X_12632_ clknet_leaf_42_clk _00082_ VGND VGND VPWR VPWR Oset\[3\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_17 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12563_ _06252_ VGND VGND VPWR VPWR _00469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11514_ _04973_ _05158_ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__nor2_1
X_12494_ _01527_ _05134_ VGND VGND VPWR VPWR _06213_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11445_ _04855_ Qset\[2\]\[14\] VGND VGND VPWR VPWR _05346_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11376_ _05274_ _05277_ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10327_ _04232_ _04222_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__nand2_1
X_10258_ _04164_ VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__inv_2
X_10189_ _02556_ _04095_ VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__nor2_4
X_06420_ _00547_ _00554_ VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06351_ _00491_ _00492_ VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_60_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09070_ _02980_ _02960_ _02961_ VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__nand3b_1
XTAP_TAPCELL_ROW_32_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08021_ Oset\[1\]\[4\] _01332_ _02019_ VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09972_ _02784_ _03876_ VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__nand2_1
X_08923_ _02688_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__clkbuf_4
X_08854_ _02580_ Oset\[0\]\[2\] VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07805_ _01855_ _01858_ _01612_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__mux2_2
X_08785_ _02624_ _02182_ VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__nor2_1
X_07736_ _01691_ result_reg_and\[8\] VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_68_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07667_ _01724_ _01635_ _01725_ _01726_ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__a31o_1
X_06618_ _00724_ _00725_ _00750_ VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__o21a_1
X_07598_ _01581_ result_reg_add\[2\] VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_80_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09406_ _03248_ _03247_ _03315_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__a21oi_2
X_06549_ R3\[0\] _00665_ _00683_ VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__o21a_1
X_09337_ _03241_ _03238_ VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_33_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09268_ _03052_ _03145_ VGND VGND VPWR VPWR _03179_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08219_ _02145_ _02149_ VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__nand2_1
X_09199_ _03106_ VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11230_ _05131_ _04876_ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_91_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11161_ _03652_ _03145_ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__nand2_1
X_10112_ _04017_ _04016_ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11092_ _04494_ _04957_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__nand2_1
X_10043_ _03909_ _03949_ VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_42_Left_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11994_ _04058_ _00590_ VGND VGND VPWR VPWR _05832_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10945_ _04847_ _00582_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__and2_1
X_10876_ _04759_ _04760_ _04779_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_100_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_51_Left_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12615_ clknet_leaf_39_clk _00065_ VGND VGND VPWR VPWR Qset\[2\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12546_ _00953_ Qset\[3\]\[9\] _06234_ VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__mux2_1
X_12477_ _06190_ _06123_ VGND VGND VPWR VPWR _06203_ sky130_fd_sc_hd__nand2_1
XANTENNA_4 _00564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11428_ _05326_ _05328_ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__nand2_2
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11359_ _05260_ _05093_ VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_60_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08570_ _02470_ _02486_ VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07521_ _01579_ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_65_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07452_ net7 _01187_ _01254_ _01521_ VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06403_ _00537_ VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07383_ _01456_ VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__clkbuf_1
X_09122_ _03024_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__buf_2
X_06334_ _00470_ _00475_ _00476_ next_PC\[0\] _00478_ VGND VGND VPWR VPWR _00014_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09053_ H\[3\]\[3\] _02836_ _02837_ _02964_ VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__a211o_1
XFILLER_0_32_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08004_ _02014_ VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09955_ _02787_ _03861_ VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__nand2_1
X_08906_ _02812_ _02818_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__nand2_1
X_09886_ _03792_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__buf_4
X_08837_ _02653_ _02750_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__nor2_1
X_08768_ _02681_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__inv_2
X_07719_ _01666_ _00551_ _01776_ _01589_ VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__o2bb2a_1
X_08699_ _02586_ _02155_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__nor2_1
X_10730_ _04634_ _04434_ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10661_ _04358_ _04355_ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__nand2_1
X_12400_ _06113_ _06140_ VGND VGND VPWR VPWR _06141_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10592_ _04468_ _04470_ _04496_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__nand3_1
XFILLER_0_23_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12331_ _06085_ _01532_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12262_ _06033_ _00899_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11213_ _05054_ _05115_ _00820_ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__nand3_1
Xoutput41 net41 VGND VGND VPWR VPWR data_address[3] sky130_fd_sc_hd__buf_1
X_12193_ _05960_ _05989_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__nand2_1
Xoutput52 net52 VGND VGND VPWR VPWR data_out[13] sky130_fd_sc_hd__buf_1
XFILLER_0_31_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11144_ _05044_ _05046_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__xnor2_1
Xoutput63 net63 VGND VGND VPWR VPWR data_out[9] sky130_fd_sc_hd__buf_1
Xoutput74 net74 VGND VGND VPWR VPWR instruction_address[9] sky130_fd_sc_hd__buf_1
X_11075_ _04309_ _04975_ _04977_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__or3_1
X_10026_ _03927_ _03932_ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__or2_1
X_11977_ _05805_ _05817_ _05755_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10928_ _04283_ H\[0\]\[12\] VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10859_ _04110_ _03685_ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12529_ _06235_ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06952_ _00650_ _01072_ VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__nor2_1
X_09740_ _02556_ _03647_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__or2_1
.ends

